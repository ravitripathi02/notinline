<svg width="359" height="279" viewBox="0 0 359 279" fill="none" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink">
<rect width="359" height="279" fill="url(#pattern0)"/>
<defs>
<pattern id="pattern0" patternContentUnits="objectBoundingBox" width="1" height="1">
<use xlink:href="#image0_1_370" transform="matrix(0.0009524 0 0 0.00122549 -0.0828691 0)"/>
</pattern>
<image id="image0_1_370" width="1224" height="816" xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAABMgAAAMwCAYAAADVqFz1AAAgAElEQVR4Aey96bOd2Xlf9575zhPGnsnmPDQpkZEcliIpUhIPsmxFsaKUbJf/zlTyIV9S/pJUpVyWHSmSODSbRA8YGw3g3jNmrWefFwApsjS4BwD6vehz32mP66DAuovPfnbX5QiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBEAiBT5nAgP785AiBEAiBEHg2CQyfzWFlVCEQAiEQAiEQAiEQAiEQAiEQAiEQAiEQAiEQAiEQAiEQAiEQAiEQAiEQAiEQAi8IAWMTEp/wgnyZmUYIhMALSCD/Qr+AX2qmFAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIhEAIh8IsJDH7x4zwNgRAIgRAIgRAIgRAIgRAIgRB4QuCX7W+27gaDQbfZbJ4UzVUIhEAIhMBzR2D03I04Aw6BEAiBEAiBEAiBEAiBEAiBT53AL4stiBj71L+KdBgCIRACnwCBCLJPAGqaDIEQCIEQCIEQCIEQCIEQeNEI9IJszcSUYv2956c/v0SYDfvyLxqXzCcEQiAEXgwC4xdjGplFCIRACIRACIRACIRACIRACPyXE2C55OBvWC7ZG7CnjVf/rB/A0+985hpMz325/uyzHCEQAiEQAs8AgQiyZ+BLyBBCIARCIARCIARCIARCIASeDQJP5FjlHHtKZBk59jOH7xBhfW6yPhfZ4zI/K8metPTk6nHRXIRACIRACHzWBH72H+3PejTpPwRCIARCIARCIARCIARCIAQ+PQI///vQU/KqF1+1NpJy660Q69dWDtej8Xizv3/QLZfL4aNHj4ab9coyK8qizqiy4fIXHzb+83173z/rx+H56c8vbi1PQyAEQiAE/osJJILsvxhhGgiBEAiBEAiBEAiBEAiBEHhuCPy8guoeJwfbhog9HSmGxxoMB5PZbLC3d9DNZrPRZDadjMfjwWq1WnCe7+7su4vlAEE2fvjw4ebi/OHq/v173WpxARI9WGvvr3X7RIb16HpB5vlpKdZf9+VyDoEQCIEQ+AQI9P9OfwJNp8kQCIEQCIEQCIEQCIEQCIEQeMYI9L8BqZ3qUGL5qcNNzMYYL0TYzuDw8Hh9eHi4nu3sbXBgw8VisbMedLvIsSFLMec8m6/X3Xo0otpmsB4Oh5vJaLhRkN2+8/5wfnE+7CiL7up7XdC+5mxZvf3SH09LuirEANf9IJ8WZk9f/9LW8iIEQiAEQuBvJtD/Q/03l0yJEAiBEAiBEAiBEAiBEAiBEHjmCfQe6a9JpscjR2zV9Wbj2fKDbjCedru7+3t7+/v7s9nuHtFiE4TXGik2X27WVBnscH8w6ga7q26jSFsu16tzFlQ+RJDd5/6j9Xq9GU9GM847RJdNeDZBps1Wy/WUzP/k6d88ZDnm3eV6fZf2HlW+s/V6ZL3FxcXa+w0NrtdLPmtWaC7wa9yvlgqyEaMdbHhDu3yGWzn2s/N0btUuhXKEQAiEQAj87QlEkP3tWaVkCIRACIRACIRACIRACITAM0/gbxJk9Z7fg4ZDIsXGo8nO+PDoZHR2dnmAAJuSRcwIsT2CyPbwUCeIqkuDYXeMdOLZYHe4GcwQXJPBaGgk2A0a+QHvblD3oWKKMsSa8YaYM+4n3dB2ut2RBq7rpsi08YpGOS8wYBTZjLvVmtEM56v14hEVz2nhfDwanCPTHrKS8+GD+/cefnj3bvfonNfbJZtceNgTH+LaqMhHW5aoMiDkCIEQCIG/K4HkIPu7Ekv5EAiBEAiBEAiBEAiBEAiBZ5jAz0ZUPRloibFusrvX7e4cDFg2OZ1MZgfT6fSgGw0ny9WGNYzGZ63HyKrZcDg46rrR10hR9ms8+zwxZrMNefqJJjOybIoJu08E2p/a23A0mvBh2eVqOBoM71L+/W40eDBGgnHtEEab1Wof8fX6arX+MvcvLxfLyZDE/9vlmiNNGc9Zgrl5QLlbrMx8l/u3u8Ho7f3D0x/v7h9+QJ6ztcs3yXXGVgCu0qy2lX29IPOZ7eQIgRAIgRD4OxKIIPs7AkvxEAiBEAiBEAiBEAiBEAiB54KA0kgr5tlPN53tDj735peG+LDJck0k2HK9g1BSTk1ZmTjlfID8OuJ8xtLKV4jy+hVq/ppiiwa4HS15V1Fbm8HQaK8d3uHBRh/Q/C7vRiySfJc2/orVmze4dxvLE5zVFdZHXkW6fYHos6/z7A1k3D4RYgMMmVFnI9ZXmtcMubU55/1t2nyX27dp68ebzfptitw4Oj69cXRyfPPi0fmdW7c+ePDg/ofnrKfEkpUoo5qHsqzyldWceeDLpwtYKEcIhEAIhMDPEej/0fy5x7kNgRAIgRAIgRAIgRAIgRAIgeeegLnC/J1nOJ7sDi9ffakbjaeDnf2DnVE3nCGmXAm5QFQpxojuWn2Fsl/k/EXOb/D+VSTVJa4nlKm8YFzXQXnP94lCu8X5nNsJUkvJdQ859iO6fJs8ZAsSiF3h2aujbnSZcoeL9eKQcvvL+cUOEq5yjPGetmt5JkUMACMJGcn8KWc02flw1D0g+dgdrr8/mUz+lHb/82Jx8Tb137l79+6t+/fu0o2irfKcMd+183aAijEkHQtDt46sDy/rfxHs7ymXIwRCIAT+QRPo/138Bw0hkw+BEAiBEAiBEAiBEAiBEHjuCfi7zRCJZESYYuhndoqczg666y+/arqvbrKz2yHITikzRpDNkV1KrF9HjP0W52/x/Iucr3AuKYaIMm3Yhs+QMhvlGJ8RfRlW5nU3HY+7yYR0YsaAIcmGwzFRZWsjzk75XMVWDSxLf+vlarEgxf6Q9saIN15vNtuzcsvcZWXfbLcbkKwfgTYZubnm4EPa+H8RZH/Gq7e5/jHP3j4/P//Jzfffu/3hvXv3GDKRba7rFIFHNUUAW+Upc/1lveh/EYwga5TyMwRCIAT8fxZyhEAIhEAIhEAIhEAIhEAIhMDzQaA3O4z2qct+7Px+Q7xVvanljdvnw4rUOp8vut29/WaINp0C7CqC6DLS68tYqe+NhsN/xFLHLyOuLvGsxJRiTEHlLpREaZGA39z+A3rhJzqOhGWkMGs7R1LEHSftfQebdrhaLk+5P+L1wPZWvOMZhVeD+cU5z4xKsx8kGOqsosd4R5263vDOOVK95oFEm9HOGWN6nb6+zkaZ3yZo7du7u7tvMq/jk7MzCy7ni8VHpQirVtFg0EOcHCFm9LZ9/EtOCrXWa52t0rr/JeXzOARCIAReDAL5p+7F+B4zixAIgRAIgRAIgRAIgRD4h0HA32C2iodLpM/jPGMuJdyGTVXUlPmWSbTf7WC0dvf29qcHRydcHI1QUtfHg9GbiK+rhHW5y+R1BNjXUF5foYETZRYyChs2MGpsxKdEGPnDSo5RHmlUgyAgjBCvVSXGN/Kr3m9WayPZ2u9aRoAhrRRt1KoIN1+5JNLDOiPju7aTwmTVc8qvKWf/ayLGnJftq+Uqco1nRKxNuul0bBvvuvSSiLP/wPM/n8/nP3jvxo2ffPD+ezepdx/Bdr5xpWUdlZ9MQLa55dXeNJT99fbM+Ouo6f7cu9yGQAiEwAtEoP3r+wJNKFMJgRAIgRAIgRAIgRAIgRB4sQkomNhB0knyY60IM3KMHSCxQINxhwjrdvZ2vzgcjL+BOHoNaXSNJY9nvD/aDAf7CKXT4WB0hgjbRzu1XSsHo33viRNzGWVHBBanSqCPd6L0mEgxlkgSO8YySnQWazVZKlkCS8k1wH+tVm5C6fXKwQ3Z8VJhplpqYWiMF99lnrI2eN45F9olvos9LRFw7mxZ17g/D67tY8M2md18tWxxayP8Fv0pyBzTzs5ON55OPmKeH8wm0/fo7x3q/JCloX/6zo/e/o8f3r/756vl4sHWh9n3mB8aM1rpHVlJRR79/NG///nnuQ+BEAiBF4tA/cP8Yk0pswmBEAiBEAiBEAiBEAiBEHiBCWhyFGKKJ/KMKXB85NrH4embX/zy1d29gy+SNuybj+YXX0dovcbLa5Q4RUadkOFrViJqQBMcCiIl1ZrkYT7nJxtLIrhwWIoqI7XqMxk1gUU9osuqLoKsa4n2F91muaINcvIbZWawWMsdhiKrXSUN/6r2VpzxXtWn7XvtuT8wYHW5oR/H5fsqQ5OWI5OYUo1mCCcbjdY8G7DEcjJgnafv93cPHN9H0+n0Xcr9f0i0/8B2l//3j370g//04Z3bb9M4Oco8GGeDaOfKMnuo5/x46oggewpGLkMgBF5gAhFkL/CXm6mFQAiEQAiEQAiEQAiEwAtIQIsz5aMguyipM0AMHR6/dO3aS78zne3+LtLqW/P50l0j95BGu0irPeK4xuWqiL4yMky91gQUpTiWy0UJKJ4ZsaWUGhihpRyryDElGs9LgHFtG157NnKs7reCbE1u/iF59m2ftzbPCD0UY+2q9f1EPrV7BsX4mhBrgs5avuv7JSqOtZddRZYRycaaSwVcN5pOdwaO1bIIM7oaLmY7k4fM/w6fP6fMv7979/b/8aMf/ej/uXj04CND5JBkRpJZ3+i7OoTajja2/hfGJ8/79zmHQAiEwItFoP3fJi/WnDKbEAiBEAiBEAiBEAiBEAiBF4uAv7e4lFJfo7khhGuIeRpMJ7t7V69evf6ts8tXfhdf9S+InvrnSKI3eXeK2Dqg7Iz7CuNiH0oWRm6W3C/RV6QBawdCrfwPEopX7TAai6vHcsrFiJgzkuwrvDgvFGREjimaKMeayyo7HLOrZVXkJ282/iEKjA0A6r3XvlaWed2m43kbLcaVB6XrbFnlm4fliW+j4HrIcDRp5kfTuNmVyzhXzNkIOOa2nvBshyT+J8zvc+yheWm2s7P/6muvTxBp83v37pwzhLn1+Nj7mFE0e+fg/K81XOf8CIEQCIEXnUAE2Yv+DWd+IRACIRACIRACIRACIfD8E1Dc+LsLdklBNux2dve7a9df+taly1f+YDyd/clmPfgnPH9rOJmcDI36Yomikqv/kEcfv+WCylpKSZjYknxgKxJ9seiyWmXlIk7LaDGjuIjMKmpr/BHyiKWUF92cz2q9JNoMr2Q0GdFhtQMlu01yW55sq7W4ph1uyL+v2Xosx+il1JPjMJdZ26GyRYjZoRJOGcfIq56FGXrJMZdntubamMgrpoGrAvPl3KY56udgMp5WLrXFYm4E3JCyCsNXEYhvHB4d7B2dnN4/Pz//gN00aaxkWOU3owEG4ALT9oeebTRHCIRACLzwBCLIXvivOBMMgRAIgRAIgRAIgRAIgeeWgL+vYIoqWsyIsfVgODohYuzNl156+XuD0eSfYcD+BWnuf4ck/FcRQLvk4jLcaj4ajtyFsg6XJyLHNF5EXtWulCOEUR99pSQbjobjwWTallQa+6VY8yDorHKOIZYe5xszoks5ZaL+FW23SLBSV60OIouada3oGmLJWBqJqHIJJM8VXvxhcCXDquDP/ShRZitVVu1FWT7qtXpWfVipIsxs1az+fDr84HioDOR+SYqylRFysJny4IRnb5Bv7XQ8noyvXLnSTabT5b07d89ZBLrAELo7gQPX6zUA23nYU44QCIEQeJEJRJC9yN9u5hYCIRACIRACIRACIRACzzcBfl8pU1VRY8dHp3ssEfzt/cOjP1muNn/EssHfJlLqc8ixMQKIkhQvj2RcVYWAESW26ZY6H6K1XEK5QHQpuAwbU5z1Symnsxn5xtwVksT8tGOU2HrFSs5tuQ1CzPsK2DLKi0WbmiTFle3QUUV/GRVmEBbrH1t0V5XBNRGJhqyqYC3S6bsMs11vRVxFrCm9XPFoyyXEOG2j4OyHqdlaCTL7dM7YN4xYS+jvvIiKQ+TNHZcDqBqUGyDJSni5Z+ZkMjohv9rLCLGXDg4O9l5+5bX7Dx88+GA+n1fb9M/yTDKduW40RwiEQAj8AyEQQfYP5IvONEMgBEIgBEIgBEIgBELg+SMwbLapG+5+7o3Pv3n5yrX/YTAa/wGBUr+H/fn6eDw9RIqNkVxzorMWnKlQkWIjHFNFiF0sFgOWRQ6I9hoYBdYvV9yGR5XgkotuymdKKOUTub583OQXcsrdJVVGTcSxBFM59dSxdVEINIdMe7TBz2q3HijMaEM55lGCTGFm28o93yHDmE09Q161avzsI8Z6KWY5n3lPq1XPe4++LLc4uzXNurklag5hxmdJbjJKDWZEtV3h/lUi8i7Bbvbqa69tZtPJg5s3P2D96AYz6ESqzR5L66B6yY8QCIEQePEI/Oy/6i/e/DKjEAiBEAiBEAiBEAiBEAiBZ4LAL/YsSJpfMjrLD1kCuDP76le+8ev7B4f/brnp/s1kMv3uejM4Q+pQgGgq6w+Gm5EKCN+kIFMSPTp/VDm+lkR9KZJcCqn0cg2isV/2agWFWR1GmPHenGL+8bCe743iapFcI2QWSyWNNCNyy2ti10pQTVjBaISYDduuwstxcOJ4Iq9KvPHcbt0yQGFmbJjlFF91zbxLpPHMNhRzPve9EWIViWa96sd2iGzjfQmzEnv2a8et/xXvEWPufIlfHBI8V/tg8n6wSzTZFaLJ3sCjvX56drZ/eHjw8PbtW3fN8l+TacLxiRyzWT85QiAEQuAFIxBB9oJ9oZlOCIRACIRACIRACIRACDybBHqr0lxLEzh/baRaMX5H0TQNyQk2u/TNb3zre4Px5I+X6/UfDUeTL+BtdhFB5NQaX5SAquAoMuKTW4wlhuQYY0nldhml71126D0bPGLPWv4ue33cPyLJch4lo7iudrmvpZi8LxGlvOJ6xAYAiiqtlUFe5aEoW6JrK498z1aRTXht69t+a0c9x8EPI8d8Vv1Rtx+Hz+qjFgOF5fsItb58jYHn/bkGY7MIPsu4tNR3LK2sdom0axFl8qpAO3YYoFkE35Tyl2H6xnx+cfno8GD/0qVLmxs/ffcRau4BRR5HktmudfyRIwRCIAReNAIRZC/aN5r5hEAIhEAIhEAIhEAIhMAzSUDNU2qoRrd1SY9H+uTelPajbn//+Oir33jrN4jW+ncETf1LkuhfYX0g5ZFGJApTGyGw2I1yrWJS/pTQMseYUsgcYhvFWJ9vjHOJqCFjKNvUlik2OdUivkoAbd/zZCupWiQZvZWs2gaX1Vzsk04ZEX0v25JMRZz5zjz6tm33iQyrVwi1FhFGQv0SWbXMUglHDrSi5DAVUvxnfjJ35fTaNm3d+lthVfUnI6LaLEdEm8c2SX9d+0MH6HiXsEHebabTWY0Jj8a6y6VtzIbj4VVafvPo8PDK6cnp8ubNW7eJPrtfHVcLtQr1cZu5CIEQCIEXiUAE2Yv0bWYuIRACIRACIRACIRACIfCcEGhCbBsdNWCLx66bEPNE7qvhem//YPzWt7/zXVYC/vFivvwD5M3pogmuj1hSiedZj/VGPDfirOSY4qgix5RARpCRcF4hZBSYZ4VSOZ5tKJbCyKOXTP2ZRisarH9vux5qqRJeCjraau22JP71ruKsthLOyVlnW9fy/XW14T1j6svU+JRjPDdizGkZkWZZttcskVURajXdJseq8vZHK++STyLS0ItNuhFUR/2+XyWX7VuWZ+5RMGRppTSMxpvziufrGRM9Xa7WbxwfHe9fvnJ5+c47P/mIwd6jvkWFIfMG5elB5DoEQiAEnnMCEWTP+ReY4YdACIRACIRACIRACITA80RASfP4eHLN7yXDKZ/50fFJ97VvvHWNCKh/tVjO/wBB9NKC6Kw+hxa6yBRc9XuM8sdIKRPaLy7mnRFm5M4iaozcYYSdKZ7ISIZsUg+1fFwDIrHIxFWyyHEY/eX7Mc96OVYyindGZFX+McZpzjG1kJtDtrabDDNijSGgjpBlHCullBflkizf5tuLKs2UcszcaZYzessapAhredI4K7qoWMs5lV3eu8umcgupVWfbtU2fec1QKWekGeWZy8T8aIzZ8VuuLb10Cm08QiQ6bDOb7SDIRgMS9I+Wi2WRotQOkWyvHR8dnh0dHa+JJLtL2bsMSg1Y02PorSHnmiMEQiAEXgAC9T8sL8A8MoUQCIEQCIEQCIEQCIEQCIHniMBW8BDYhc0hdT6fi929/e5bv/Kdo4uLxe8RofU/8+7bCCgixDbnOCAjl4gyW7OhZJNDJcDwNUZzbRBLfhROLq/0qGWRdcUPJZLXmCSF02NhxVNlETFbPyOzevFU9bb9WacXb+u1yf+VZK0DE+V7/CJ71Pfl+94q9eX6Grbz9Hy8dl6+91oJ6KH0qg0CtuKsH6dz8kOusZJmPleuuWTTo0myJhN9Z0Qd7RKwhgbEDJq4n2PBswVjGS8W8ymRZK8jLA8RZY/effe99yijJLM1ZGZdtDA4O8gRAiEQAs85gQiy5/wLzPBDIARCIARCIARCIARC4PkgoKgpufL0cJVjEyPHWFbZfftXv3u0XK7/kB0n/zXu6TvL5WoXpUOwFXFXm80QIUUjLRqqPz8WVFzUTpUllsippdQyOqz8kDqKvvlPEVbCaqMQo3UKlHAyWow6xKrZA38s77LE1l/fT+u3iaYWvWbbfCjrp5+lk+yllNdKrrqn7OOdM6uMb1tZ+1/bH00ZBWd5Nieo3S6XS5Ltr5oM1Ck6tybFWlRZk2Msr5wYceYzcpux3NJpeG+EnHN1R0uH6r0XROl1JOcvdkMFGw3BsbYgQIi5I+j145Pj0cnp2c1bN2+9S661Zh+7AfaOhpz73+royfxty/+tGk2hEAiBEPjYCESQfWwo01AIhEAIhEAIhEAIhEAIhMAvJ6BM8ShBoi3xdxHN0nw8mXW/+t1fu7xYrP45EWP/Binzm1iiQxURZbRjljXajFOTTQonPxU9RlJ8ZFrJn9qt0nLuWmnhvtv+AvtU7SCi6jVl272LLZsMa8/7iDKf+aGp6l85tq1j84g1I9AqEI766DZHTG9NYtlWq9/qtbbboPrnPvOwXeWYZ5d31jN+WE5Ua6RZOxiPfbk2lIMVkly3CLImyhxTG7/Sq545MtpUzslMUdgkYmvfluiFahxYQdjOKUoI2nA8X8zP9vf2h+Qku/vTd9/9KX4Th78AACAASURBVC/Pq3TXEUnmiEH3Nx5trNt6f2PpFAiBEAiBT5tABNmnTTz9hUAIhEAIhEAIhEAIhMA/IAJNKjnhJnm2U/f3kIoc29nd7775rV99ibzx/wvi5t9R6rvImUNzciGfcEMoHV66pNGYMEWYSfjXSwQZYqyJMpLyG3FFmcrv5U6SHPZdye5pq+wPgshoqia0LLGVTOWiiCyzTv3kjVX4oXiqp1y3+yZ6hsNxlSHBfeuHe9QSSxrZb4B+uajzkHt1GesYa7wlpezIp1tn1ERXuxlT3jHTUu1IWXOg3Wqbs2JMyVX3VBkSKVasHHm1a7cKsybIzKvmx4gyxd10PC0xJq9awkmoHp1Rh7a30tF50rurL113yQrM8R6nq3v7exenZ2d/8cHNmzfXtWunSy1ry07KNU7O6xcf28n+0ve/uFaehkAIhMCnRcB/xXKEQAiEQAiEQAiEQAiEQAiEwMdOQFGjbHnq8PcPP0QcDRfD0UQ59irl/kfE17/l+W9QfsfAMJ4ZxTRakhsLI0Q7RIktFiXCSooRBbVC7qxWPjM5P3KMvowgK8Hz1/suceRYHJcfD0WS0oqnda/gaWNukmn78LFwsmiL0nqS6+tJ3q/2TNlku02etT7MBzYek2DfP+Y8K/HWxmIf9mmd/nDZZ42L/vpE/fbbH62NFhFm3dpEgJf93Puynvv52o7LQvux2ZbzKTFW15WXzPfEjY3pfsir1ZJ6o5KWy/X+/v7Bo6OT43ff++C9OxvXaxa3zdYKar9+5vu2i+3xhG//JOcQCIEQeJYIPPkX9lkaVcYSAiEQAiEQAiEQAiEQAiHwXBNQyjTR9DPTGBPXZOb4xXS2x26V33qdSKw/IRn8v0GWvYXnmSiXPBYlw1YammrHHFx4s20uL65Kjhk5piRrEWP2R0xZKRp1jGOo9P9KnJJSTVw1YaQoeiKqKhCqlmq2ZPtN9Ch7WqQXTW+PavnJ3LaRU33kmWMk8z3dtQguorAqEmyMDFRG7bAb5XQ6aQn0fcDhnPtdLW3HKDfzqTlsry2m1PLTyzLrGQWmPKy+GB/ar6LFGFwxkId+sdonfxmRYPXeNoxoa+21XwkVd0uYlo+kbcVafdBkfBcDuiKF2eCEEi8dHux3Z2dnP7x1586Hq8XcnneoQk+KzwLVJuYgHx8+r3ePn+QiBEIgBJ4lAhFkz9K3kbGEQAiEQAiEQAiEQAiEwItJwN87lCZomjFrJUeDb3/ru2+y/PAPl6vVv0bUfJfXyLHBnEilDUsoR+xEaVL+qtZ2jEQ9VZQYFsalgJuf20XSZ7UMs8kp5Y4CyLxbXlfie4SRzzyUToqyNqxtm7ShbOvF3s+eW9RZ/6wa4YfizGeKLc9NTfli64gsYF+8sb+JSzJrSWN77zPHpBDzelurXXNv5Fw72hvnYrmSV1uJ1fpv8ylpRgVzj8nJcfjePvq+qp+eC+3blpFlFCxx5tJVyyDSHJDAWEI5BM2a9ZnddYTmyXQyeXh6evrjD27d+mitveRghHzPJcHqh89yhEAIhMDzQiCC7Hn5pjLOEAiBEAiBEAiBEAiBEHhOCSBb/L0DQzNZj8c73Te+9StfHg4n/5Zllf8aSfZ15AxCbFm5xebzcyKW5sMlisXcWsaDlbApf8MySyROxYghcUpIVfSYPqYJqCaCFEItAmpABFZzVUofJVITReizWpbYizPbKqFk6yWlmliiJVvmD5KNbowOs6yHEqmVrcFtn/uM0Sin6rB2O9wRk4T33fn8vLvgvDAqjjkiCast29vas7a8kmqMuj2j0ZrvVl451hEbgBoVNiGvmMs57dd5I7A6dpssV9XPq7XdRiKjko89Qypar9hVwn+WWrpjJn1MpzPDydpkDVWDBkLtjGG/RDTc5sqly395987dRzgyuyeSzBPDhpuVahBt+vkZAiEQAs80gQiyZ/rryeBCIARCIARCIARCIARC4Lkm0IyMEUjdZM0avRk5x748Gk//p9Vy+SfM7JvYlBFL+C6cJZJsjHAaKssGShmOXgq1pZZrIqMUL006Ge1lByV/tmfWcHZj6rqE0MioWk6Ip3E5pUcvzkxcP54gyzBkK0SRSzE990JHzWO7vVCjOH1736K3zA/m2JhTO1OzH4eiyePx2ClndFtJwG3ONMdekXAuk9yW9Wxdx2371R5nD3/aXj++btP6tQ2f9/OcTNj7gMM2+mg42/Haw/e21Y+RTur5YynIneUVd2pB348nE3cSpcoQZ2besW7G9StslHA0m04/Ort09sP33nvvnHdEktkgg2sNM2DHnCMEQiAEnn0CEWTP/neUEYZACIRACIRACIRACITAc0RAOaR0KTHS7AvRRLPp7vib3/z2d0j+/idEG/3RaDz+MiVct+fcKs8VsmeoWnF5YKtv1NR22WOVQn4hkKp1pJBiaEhUFun8S3QplczZ5eFujZazLWXQEBFmANSI3RxLnG0jpRRnqC4ivhRWjKXPKcb5iRxTphGtRVt+FEiKMT/e1+EzPo6pl1/2b5s+cx7KLMKyuo0fe0VC+e7pY2Q7PKgx074RbI5Dv1f9bvtw5WNft5dk1rHvNiZzlhn11vj5TEFXY6CNCXnIfLZiqaoxeUaMWdZxeRiZZvvL1bz6ZrKWx5KNkGXdcAwf2J0xruuz2U53dunSD27duv0If8aEBju2wocJP5mf488RAiEQAs8qgQiyZ/WbybhCIARCIARCIARCIARC4LkkUBIES9UWNqp6ppOdo7fe+va3uf5DEsH/K6b1FSTZECFzYc6sFjmmGkOqYFx68dNHPZVnQbcos9YVedXyj2F7SvjY47CElpLKRPYtCf6IZPj98XREFhs0Iojar0LaHqPTjJhyKaciqPVvf8qpbcQYMsl7I7A8K5d6IWYf1nky3nbvsybejPJqkWJcVD1+bPvpR7g9896jZ8AS1OpPQWafCq4SZVtB1o/x6f69loNnhaFlnKP15NezmExob9ufX1fNB86tPkyViNt5jhFmCEH85pjccNpEtgtVhA0Gr5Mb7nhnZ/fB4dHhj99/7/1HdLPEWzoRRl3f6xNLVrPLjxAIgRB49ghEkD1730lGFAIhEAIhEAIhEAIhEALPMAE9lkrq551He46CUbE4fgoNu929g4OvfPWr3yHn2L9arFe/z3LKLywXCyXLZrWcK5VwVGuFGmIGUYWocUdHRRVhYdVTSS/vaXu1IOIJ2dMLnxJDyh/qW25nZ6fb3d3vxuwW6RC2+eNrROYjmyLHxpxpGnnEsk5WDC7I13V+cdEtKoqqWipZVJNgLIojI8tqeSbnEZFZ5f9ow40DGDhnVhcageUc9EcGT9kJ/5Wg8p1suPdQeJWo4toevbYdyzYJ5q3xY0g5JNnO1PRelC0OT6LMeFDjc1mpAk0fta5lm0auOYb23iWlHuZBa0w2tVOoYrGXYwPWmZp3TBG5oZzuzHptPI6E50biDUcbnzM+XvJNjYZn9HV1f39vdXZ68oP333/v3F1G+b6mdukFnxwhEAIh8EwT4F/DHCEQAiEQAiEQAiEQAiEQAiHwtyWg7/DYRkK1G37W861aUeUMN+PJbO+rX/3aN1Auv3+xWPwLhMpXEWIuq5wjc0zGT3gUBcvjIF8QT0osD+VQtVnneoDQmSN/2jJBl1UqpEzk72HvOiaTyvtxKeWCJYUlsKpEi8BSjk2JLHO5pSLLBPkXF3OS5iu3FETbeXHdxmC7JYU4EzmmHKM3nymOVuQWQ/pVP0aQ9XUUeFLwMP9YHYxPyWTdvpzPvW/ia1uMew9lWTWilEJ+Gb1mrjHrtmWoPSeKUUdpZbL+im6jquUUXh4KuGqPe1t33h4UqYM1k/W+n7/LP9lsVMQ1vrazpXKRr4ywNL5oB0fato2p23Zp+w0iAad7uzs3iOD7/q1bN2mZgfNj+6l+8iMEQiAEnlUCEWTP6jeTcYVACIRACIRACIRACITAM0ngl/mOeq40UQNtZjv73Ve+9o3X8Sy/N5/P/zlRR19ZrjZjk+ITbbQZGCpmEq8SRuTKahFJVdtpt6iltiSwFz21XBFBZiSW2sXnRmoZKaWJqeWEW8G2IKKrz/+lGPIznU67ndkUyUTuLUTRgmi0+XxBRJWizHZspR1NWrXllQqnyQg5xdk+7U+x5FlBpgCzrs+e7tOyBk+1c82USgqrJt+asEJEOXqKlsRSlvlHNBxVhmiuXqA5Fudhmwoz72VV5awgfRgMGW/bqKDlJbNMSTQFm+X4qdBTIOrjXGppGy49VYYZLedyTBqp50WGHy6J7UUc5ZlctyFv2ojTAK676LLBzs7s4c2btz5AmJ3TDwGB27C3mmV1nh8hEAIh8MwRiCB75r6SDCgEQiAEQiAEQiAEQiAEnm0CyqNfcmB1avHg+qtf+cY+Dux7yKc/RLZ8j4ilHRzMgsgq036NWMJHDjK0SgUi6WGUTxiUfg0iHbT3yBtEjYLH5ZAuEUTCVASUUsehOB6ljYeShy0zKd80UP/MyCvF0pSE8vbqskqjpVxaOV+09u3fBp+WY7bX6s4eP+/nr09TMFX+MgVUHY7JF6q7FqXl4zaXtsTS68dt+I5PSTHlnvMxDq8GY02HhCjkU7ttOj4k1tgoOEUfMosND0pweV3GirH0kWSKLsWh/EqkWZ+PvbZxVBd4O6PSGsNiWU5LcSZLhNlW0k0mbH6wbWNMBSQYcWZyYE7DwS4/Tqg0n0wnP7h1+/bNbetZatlA5GcIhMAzTCCC7Bn+cjK0EAiBEAiBEAiBEAiBEHhOCOhIOEhi1Q3Xr7/xucP9vYO3WFb5jxFMv0W01pXKG0YIWIu+WpuDDJdiEvwWodTclMv8VEUcBjy5xE9RhJBxaaWXRn6VO1LY+Me1frQz3UZTbbxH9ChxyJLF7pMuOSQXGjm8Zrs7FXGFYSJybNk9enTRnc8vkEMtyqvWDVLfCDNOdst1W9aoGDJai85on/e06dgcSx811gsn+64oN6bRZBRn3NOYH62MwquJsQpaszPb0o/ZbrutARSX4lS3CDGfdN1stssYxuRb26sIuIqikxPczOHGYkv6rhRhJc2EStgez9SDjlt2PHs8d8oiIm3dMfZ+0ZnIwXkoAt3dsuVLa89Kvm3YCpOvhiLuinAMm4dEov1wPr94++HDRwvq9jNqg6dQjhAIgRB41ghEkD1r30jGEwIhEAIhEAIhEAIhEALPH4ExQ+YzWO3u7XdXrl17aTlf/lOiwf4ZUuVLSK2x8oVoI0OUlGO4myaxqMMjDUyLIFN2Kb2MgFKS+UqZpsgpqab0cZkiH0VPn1urcoNRd4TcUvAoozwUZ37YZRFZhr+hn4vlonvw8Lybk6NsTSSZcVc1HrvD5TgGPwqxFoFlFBbjYVxGoRlR5lHSiPEtGVs5rm2usU1t8KiEsl3EEmdGVfdOqOoxxvJG1ZJTfXJfEm1bri/j2U8tfaQ/I+CeHudkKn5ZtQYVYBVhpyxkDOZeK8HF/D1btyrIkPcbl5halR9yHVGuIta2LJrYa3NWvzkOx9MYDf1uB+hPcv4TCwgrThe7uzv37t29e2uxxEK2HQuedNqGmZ8hEAIh8MwQiCB7Zr6KDCQEQiAEQiAEQiAEQiAEngcCv9Bx8FBF1K1eeeVVI6zewtP8ITmufoucVbucWc1YRshllbgoiivE6qzUIioJoVM5vkrTNElVNKzGH5cyomSQO4tt1FMzQUZJKWR6WaTcmSBvPKaTHaTYiCir3W5GBJkSzJxjF5V7bM6ulctatlk9UGdM3i5Fk9Fho6H5vcYlw2bsiGlvyqA+isy2FErKL8UdPxidEozWeOY9L1FJSCTI+LwjgqsdPEAuIZRKXvmsCSspMnc+/EcZ/2ssfK+YGzAGhZfrVPs8axX5RlTcdDLrhkS6GWXGAlKGUD+b2ONdcWQ5aSkw26BN9kqoqDzbd4wl9ShhXdulUD0v4Vhz8LvblHDsmSvK/F6pZnt+v7sotGOk5cPj0+O/eP+D9+61+W80i5brQVglRwiEQAg8EwQiyJ6JryGDCIEQCIEQCIEQCIEQCIHnhUB5EAZb8Ub9DcJjsDq7dGV0eHzyeXzYf48S+8eIk5dNgI9AWg1YmkfkEptHUkUBpOzhbCSS8sQIMM/DcYveUr54KGxKQBGBRrt1T7RS9W+ZPoLJvFkV0VRtNpnk8kiT8u+Qd8zcY4q4c3asfHh+XnLM3SeNTOvbMcLMyCnCoKpdhZTtO1PHWQdnyzsm6zdBxniIGtsQQVZyrLGhnDYICcaYavXpth3nVMsgq8323rlXudZL/Wx8FGaNRd1vJZ28FGkKQcdCqaozYs7THXbxtG0e2W61vY36Um6tiRarRHDKr62rsi35OrdWB9nF/M33RkdltdqgGmcdoMc2mo6hDQaMAyWoGexm5Ce7hmB7hNj8s4uLix88evgAGBtzkYkzggwIOUIgBJ4tAhFkz9b3kdGEQAiEQAiEQAiEQAiEwLNNAMGiZFHW8PH3CTTMcOOuidevv/Qyb/8piuRfjsfTryHJdjYk28LRKMUGJJfHMxGVxTLFXsQonioyijaHRDNp3PxUonjljr6F88rIJ14YSaZ5ap6NKCzdE2Mx+qsiqRBsvpwgimY7026P6LGdnR3O5OpCaH304GHlHTOXmXMw4ZdjMMeYZzcLGCrvEFFaHO+NorIPx+yyw5J2vDMJ/4rlmit2zFwh7Ryr4+6llOWsVz6IU/XXqyHL8cdnJbDkyv3Yfihby0jrvUIKEQU3j5r39rnjcUlpHVQvVEBSqE1gPCL/mmc2SGAjggVflJsZGNHW2lQ0OkaPWgZKW54dl1F0ijeZq+Hk5KGG81ty10/HvjtDKtImZsx7IgUhy5LaCWJyMp0tefxTXty4dfN9DZkmsSdQDRaTajk/QiAEQuCzJRBB9tnyT+8hEAIhEAIhEAIhEAIh8HwRaJ5El+Ph7xMapNXJ6Vm3v7//HdTKHxN19buLxfIIUaJPqnKIHAKzEDdEafnQ5ZS1XFH9ggCzWYWM0sejRYu1TrymUC2HbPtCWn4r6WjTpYJKG+XRxKT8XNeOlUoylkfa5oT+LubzkmTulLneCjeTzJuUf2zkGOde2FRkGvc1Ag0Vh6LJw3EuWaZZSxhXc+Qdif55ZzSWkqwJMqPdoFHiS1xtLk0B0khJqtZum3ObjzPxvqoxIZeQ1r0z3I6jCbX2XEE2ZHll8SRKz3fmHnNXSuu6SUG1T/dKQUojzmDPfNkzoY2Z8v3hRgEFsuq3Pts8zF3WpJjDkJVybYK4k7E50dpRu5O2L5FiCNFzxnj7o/v337m4IHSvceiXWj7puB9AziEQAiHwGRGIIPuMwKfbEAiBEAiBEAiBEAiBEHiOCTSzo+0geGg8mU5eeeW1N0gq9jtELf0ThMqrRI8pVJZbwYMnQVzxMRJJOWPVJr4q8qjEkjx6CdOUF6UUTn6qx1JQJaZcQmjbRi8pdIx4UgQZgTUmEs0oKsUNuymyxBJJVj06phb1VSKKquYHU/iwJJDOEFr80do4Ds8l+LigZi1NnCPZfGc7G6LHlotzyrj802WfVkBO8an3nB2jn4pU49xHrlWkGuOtfT8ZgBFrjKT+UM1mag5Gezn3klI1Z/jxp+1ISbu8c0mokWo1D6Sgg3b+jtPIO1nVB5lle06serICB1Ff9NfEXps0bdZoLMryVyUkAzJCzy/c+cndPx4rlmHOzN3GA77/Ad+rH/vn6xhMZrOdm9PZ5D998MEHH9bEuo27XXr00WTtLj9DIARC4DMkEEH2GcJP1yEQAiEQAiEQAiEQAiHwnBIwAkiHguAYdlevvXSJyLDfRdT8PtFLb5Gba8dsVBykHKuoLHLHTysqqhddvvRQJJkTqwmeJlzqhYaIQxlTwqnORkE1mdOWLvqeuogaI5rID18RTUaRTafKMc4lhRRVNIYwIg6MbTSRPQo1dI+fkj1KIz4qOH7ws26QP0SLbZciLkjw76F4YiCUU5qxvLLGRB9tzlWmzJVtcPSRX3XeSinlUj9nn9ufifC9riWQ1tM4be9rAjQ3JlqsIsoYrJKtLWFlHtt2XcJq9JtSTrFoPWWVDMdGpinleFfluHbHTQVYzanGy1io51JRz7VhgfKuTYVxMlKa9bDLkn+OHdZ8BkTZMWT9WC21nJB77ojK98mL9pcf3r/3w4tHD6lZcWq2uG3J1nKEQAiEwGdLIILss+Wf3kMgBEIgBEIgBEIgBELgeSRg4BVOZsTSykvd8fHJV8aj6R/z6B9fzC9OWEJZqaxQPZTZHsoZjEqLCFsS2YRsUuBgW0oWQaH0mCJnG00lmF7uGMm0eByppVxSziiTuNjW2SXXmFKM1ZzdlPNMQYYs2+FDBnnquMSQ/kimj1rqJmXEeGYb3BshxalFeTEalyouiQxzMmuWEDZRZuQY9Sm7XLK8kvcuZyypRXlbcjy1xJG7SpZPm4qkkoacnakbCHg02eV89EVNiBUP5Jciq9pjfOo8uWyFY7XXIssUXrzv+bYa9b4S6G/fKccUXk61bZRg30jFCc+Zn220FPvNWcnbwhXBJjvqC6dyw/muPo5ObqP6nur7daTD0ZqqrDpdjUDDsIdD8sHdJ0rvzgfvvXuHOprGXo7VFLnPEQIhEAKfKYEIss8UfzoPgRAIgRAIgRAIgRAIgeeKwFMyY7hGim3Iy3+FiKX/DrnyB4v1+nPLSlrfzXEiBCthqtAsTdQou9j1Ucm1XtSSvV6OuXDvifhpkgjHVFFPCh1zlil3FsoohZriZhtdZV3bn1Uuriaapi6rnLKbI2Jsl6V/Y+STyeTH1Jmg9mY895m/DLXdHFsytebHlFzm8WJ5IlJMeabMW9O3ZRVlGDYGpzRjuSXPLFPyyZo892iRVWURaa2eeNOkFFFeVHwsv5RMlndeyiYFVltC2u5N0G8bSiqXp/oluFy1hBlCynY9jBKjcp2NIvNeodWWtrZIPCWj0WrmDqvcbdVna9cQOudR7VDGs7Ku2ilp2frw3q6ejJvx2B5t1aYGvGEYYHFny5rbPo/2T06Ozt+98dOfLBfzu9bm0BI6+F6W+SxHCIRACHwmBCLIPhPs6TQEQiAEQiAEQiAEQiAEnksC/P5gKNGAvGM7m5dffu0ykUG/Q2TV76ONfmWxmO/xXnFTVgSNgiJzNaZixaT2Ls9TLiHEFCws7zNGykgphZDCR2njoWypiC30ifXqg5wy35dyacRulZZRACm+zDu2566Vs3G3byQZ73bYEGBvZ9Id7s66A95NGdbOVpgZAqfYUmgZXVXJ+vF5M9rVN5WGItKMNGr0Z8QZDw18YsyOxaWZHs5H6afn6SOzeqlUook+lF8VnVbXtuOs2/PyQzwqk2gfllHdIavk4dE2C93KMx6N3LHTcrBVDsqALUKpt23XdmRcfrJ62H5tlNBs8alNCIodSzYt539ILqPvnF8pqyrqV0l7ts531Mux9ozHDpxQNsXdkPHy1SjyQDFSjvmHvwbdlPPl6XSyPD7a/9GNGz/9EbWUYlW7Wqg+uMoRAiEQAp8RgfYv7mfUeboNgRAIgRAIgRAIgRAIgRB4rghguzAh3XB1+fK17uDg4E380h8hmf7JZrW5QtYp9EhFHBk9pPwo8eTjJpF0My0fFnFhj3WOgmboDoxKHz5GSulxPMzvpShzqaURaL6bTNuvMUqqCXWn7MpoxNj+bFrLKV1Sub+7w71ybNwdIMgogiBDptFmCTBdFBdeG2nm0kvbwY/xrLVrlBmhYyXQKlea4qgGhjQq7+MItwNt867xmYjfqK/+KFFGR85N+VVzRCY12bSNnuO9kV6+d44VUYeQsvmSYJT3OSOuZkfmIhOx7oqj5Bb1+8O2e0FW9axL/7VzpWP3vf3QrtF47uTp+4qU42z0XI2bBj37zqPGvm2ryvMXYIhtVNIp0EYsHbVdJRs7ia7Y1EARxuvhhF4nhwd79+7cvn3r/PwRSy07l1oKkKbq70sPk0c5QiAEQuDTJdD+l+XT7TO9hUAIhEAIhEAIhEAIhEAIPJ8E+P1hMDg4PFpdu34NCbL5FcTGH+BPvj2fs2HlZjDn9ca1lViVEiXKlV4ued2WSHJGoCiSNkQfDZQzCDKFi5FNyrCl0VvIF+WYn4rkgpkixratX0smud8lUmx/d0qUGJFiezvd8f6sosYOdyfIsSnvkWj4HeWXUVlKNcUXQ617o8ZmyDEFmdcUp86YfGY8p/yaJaGOQUWksKtoMLWPc/OzHZdj11g5jw1RYi2aaivGNHGVm75JJqPCNoy9Eu3bsgIKR6Qkq9xijNGzoqy12aLcuGmcLMefPrpMlvWOMVQb3CgmbbYi3mjb/Gxe+z30Sy2NVJsgtdzYoIQZAs56S2RkDctx85+zrKg1v6OSeX7FyrEm+toY4YuorHpN5NHVBpfYJk7U32w0HrHCdfLhe++99wMofSQrjiy1lEKOEAiBz5RABNlnij+dh0AIhEAIhEAIhEAIhMBzQaAshiMlQmjz2muv42Amr+BHfhPh8t8itK4QQaaw2QxacjAVClbFHRTNG+YbRVlbZqluUXCVHFHosGTQJZNGQfGqlacvdsMsMWXUGQ8RMwgjzmS2qmgwpZZRYseHO93Z0SGfve7S8UF3hCS7xPXx/k6355JKRqPsQt3Vsko7cZjmKjOqbIc2XHo5pX2F2GRsOWUaUoq+7K+kV0WwteWcWjGlUVs+SUUO59gfOsI6EFBGqsnD902eMX/kWAk13JERWFa1LUqUNCtfphwrIaU8tLW2zLFP8K8cq/Z4WSylDkNFFz+qbv/FOR7L+Glur4kyl5YqviYTdhmlf0ZSEs2+FGD9nOrMIGtpJuUpXP0oCLcja+3X9+lmAsXEHzQ/IGm/e3yuZ5xPrl29cv+992785/OL8xtVuQkyL5vl2z7MKQRCIAQ+TQJPYnA/zV7TVwiEQAiEQAiEQAiEQAiEwPNE/DVcQgAAIABJREFUQM+C2xisFSQsnbt8cXHxq4PR6LssxLu0RKSgUigwMlqonAzFKhJMWWNEWL+0UtHCLVFa5rtiaWPJsfZrieoGddQtSH6/IGJLQWbEk3m/xgiXMZKrwrLoYobYOSSv2KXTIwTZLmLsqDva391KMfKNTRgGQs7+7fPhw4fdmjglm1suh/VxXIOdJnicF8sBKTvo5st1XS8p/OHDITnNSPY/uegeIdHu3P+om6N6prNRd75g6SftzZ0fgOyrz6HmlwsvfiLGOBshpzNrzzjzfI1U7IZKKErRv/U9l4xivsonyw8JafN5seB+xRgVWh61dFUBZzn7r/dExm3nXcqLdqxfB88nRNwZOWZU3GbJ98H1ivNsNqv6U2Yjm67b6Rab87o20s3+23PGq0yjL/5rZ5LKOe72fXE2uswx8J7otjXlHSqDGB7z5vP/9fd+44v/+//2v/450vQBHdlZ+yJqkPkRAiEQAp8+ge2/kp9+x+kxBEIgBEIgBEIgBEIgBELguSHg7w3YqeH64PDY3GMvrzabf4oQcffKl5EmxFwRcYQdIhoK3UIWf2SKn16aPIlGarmqKloMgTJleR9RZyVZpGEdc41Z3h0xjeKaGl2miEHAzLjYR1RdOtnvXr5y1l05OeiuIsmuXzrtLp8YRXbYnR4ddIcss9wjkszll0aDzThPptOKJHMp5RQ5d7i/X23vkNhfAWcZc5m5zHKH5Zom/je6bA9xtM/93t5uRZ4phdaMzZlWnBTnkkUaMKUWfzBiNfcN423iqkrWtfduXqA8cp7Kq4GRZNQ3kk5T1Oo08aV0a1LLe8u4JJXy1rMtGHnUbqHcO5Zaimo7vKtyPFPU1aFQ46JEHLLPw6WcLh2tSD7GYSSZ7bjcUnelGKvy3Pm8H5/te+87njKeJvqmk1k9q904mR0yjir00OY839vduf3o0fnte/fu3ab9eXVC0w5le80pRwiEQAh8egQSQfbpsU5PIRACIRACIRACIRACIfC8EkBcYF44Dg8PER/d0Xgw/jLS44sIrRmPF5ojEsCPDcpS+Cy3QgXdhV5BJLlcUOli5Bi5sBQsJdAUMwQWKZu8J36KnGS84zxCZCle3JGSTFaVgP/4YBcBtk+02EF3csiSSuTY5dMDhNkxYosll7zfuKyTTy3pROBMkGFGhyl7HFuTPUSK8Qy3V2OxH8fETpzb90bA7dU4los1kVRd99Gj8+7K2SFRZA+692/f6W68f4sIM6ZOu64NVFZVTjHaWhG9pu4x/ZZt+8doOUs6z/WgbTjgeOy3CS0jr5RSTUKxLrFY2facUDXLKaMojPR6Mm5e8xyhyDg896LMtu2bh0ZxtT6UeraxNucanBmHZVZE6S0N8Rq43JX8azu7vEMsWn9eo66IMyPDNHvynQxJyM/7YkoEWi/KjEwbjeY1DosTcWhkYXE9f8C8N93l+Wj83W9+/Rs/ePtHP/gRf7ceOQeOPoCDWs46RwiEQAh8egT6f4A+vR7TUwiEQAiEQAiEQAiEQAiEwPNGgN8bBgPEy+qll19VdLzF8sDfR3q8ucKAcNYGoVPwK5wUJJ4VVBV/hBwxJ1XtmIjY8ahoKeVQfajNM8LQOOtGFGUIIaTNDJuygyjbY+fKS8eH3UuXDrsrnK9fPu1eIoLslauXiBpTmO1WQn7zipHgjCWGSjfarIgmYpvo36gwo6/csbFykJl3jKWKM3a/nBI5ZhL7Pc989twRk90vjUDbZUfMmXnKeLa/N+tmRKLt8m7KO3d9XLoUtJYkMk9mrIAa886cXiPzi5Upc27tnUxKdHmu8SKZ6NvD/GKKMCPPPIwyM4eZ78cm0qdN6/qnBBj3FCDarYm2XqJZRillGa89K+aMEqv6j9tpSyMt60cOvrc9xy9LB6EYUyzWmKrdNt6+fQWo13RQ41fSee/3vG2bNZbrDeyILlztEnm2t7u3e2dnd/fP3nv3xvuOm8Nk/R522q7yMwRCIAQ+JQKJIPuUQKebEAiBEAiBEAiBEAiBEHiOCRjOs2ZppfLkANHxEjrlpI+Gcl5KEA8ljNfKMUWLbqjkh6aHo3KRKXzURgqYx0fbJbIzEb5ijSWMuxiz/R0T7U+6w4O97oT+rxLBdfXSpe6I+11ykB1wVkJN+FTeLSWQ+ojuVoRAVUQAokZZU2NE5DiulVFONQbFUctV5thdVmn+MyWXM7IcMXGdedYW5CYzyurk5KK79OCku3Z2mfGcdj9572b3zo33ulv3HxLpxTwmO0jCOX0iu+y7lik6HqWf6oe5I4RcGqnoUjK2qCvHSBTXFPlGPXOUrblXTM3PL7oBsXq7+3s1jzFtO15Fn3NbkQ+teDNmz/RaYs3scP3cfW6btZQS2UYwGUqz5V5bO2fGcvFobsRXN9uZVL87O3s85Xs1IpAotovFBXd+z+4CWpc1nhHtmTMNQ1rjcsdO85rtkL+NcdJ1CTu+kgpzmzy8OH9pfmf+lZdffe3zP3n3xp/dfPeGa1YxcFtYren8DIEQCIFPjUD978Wn1ls6CoEQCIEQCIEQCIEQCIEQeJ4IqEDKj3DaXDq7skMery8gmn6Dz68jdU6MXuLQjXjBirs+IkmnxlEWBmHD0sr+sEEjiyqvFgKoRY25LNLlinx4tk+01gk5xNyJ8ux4t7t+ety9eu1Kd/3KKXJspz5GeR1QZqKEahFIj6PXFFzKqIqYQkS1aCbPRmGR5N8oMuoZTTYlkmziGcnjmIwMmxC1Vs+QVYoso8eM4DLCyrxpM87mJ5twfYi0Otw/rEg0BdejBw9LGpmTS2GkDDM6zU0GJtWHko6x+Y4Pjqv60MiVTISpY5sqyuwPYeW9QsyKtYQSaj7rn1c0mwKOvkpG2S6yz8PvxHLW853tOCaj0VwKW98Hc9yUu6KebZQuMzKNr5VySj3V1RIB6FFj4Wx7NQe4tusmPZWf9juEa0UJUs5qSlXKMZz6LpYUuXn58uUP3vnxO/cYKes9pVA21Ya4zhECIRACnw6BCLJPh3N6CYEQCIEQCIEQCIEQCIHnkYC/L2g2Nsqay5eunJB0/TtEQv0mAURfJSn/vs7G3F5IFfNMIciebEioaFG6KK8UYkoVn3k/KAeCLDESiQ/7X3a7KJE9xNQJUuxod8qyyVl3/Qwxdv1K99r1q90ZOccOkWMHCCmXPe4SXVaHUk7poxQi6qwipOjPqKZhLfUzX1cTPxW1xYwUVo5FaWW9WsLIMs5+6WdbgqmYInk/ckwhpgw72N0lWf9eXU+ou8M49hnPEZsDnB0fdyecZ8xhcXHRXVw8IupsoQlr49T+FA+XUirN3IBgTHnEHALLMTWZRl8KJ/qejBFzCLKd6Q5jYdmiHM1HxrVfjSKqZBTzV4CJ1cT5LiX1m/O8IS/ZhIiz4iN7OREV5/fmJgG1WybtemikHEPlLKO9ldt08r2wKcNW9rkLqJKs9a0EK2HHOOq7pbDzMGec7PzTf//0y/QZzXo1VD5yjyMcrA529+9evnL5nR//+B12tKwRMJj6C8KNnkx+cWVAyBECIfAJEmj/Cn6CHaTpEAiBEAiBEAiBEAiBEAiB55aAOcUwFMP18dGpYugKM/lddMVvLRbLV1hMiaVRXrRdKz0rMpQm9RARQ/364GLqMGrKw+CmJsZIBI8o2kUQ7e9OulPk2AFLJ18mUuwl8otdu3KJ3GMH3RGRYofkGdtn50mFi7LKqChb6/uoe0Zb0VIub1SAEQ1WEUxIKkVOk2KcGYflFGf985JNiJvK58UA7cd3fiyr1FFMGRU2MX8Z4mpKXrMdxmvkGTsz1i6YCrP9kmhKKmKmEErmKkMPlQij2Zr/RPnGPCRcY1bq0Y9SS4HotZLMjFxPj8M5MOkWocV1iSnmUdy3z2Uslz6KzGgxj2qzytStzdSh9JKTS0ptZzhQji1b3jPHwDPivtoyUeooO/vv2QbcnKDmUOKOB4ynfS9Gij2Wow5S9Pxt4C2BfNTaRZh9eHhw9Bd37tx+7+HDh1TekIus/sIYMmfzHNu/QO0mP0MgBELgYycQQfaxI02DIRACIRACIRACIRACIfDCEOD3BRQSUT7Xrl5XxLxCJNk/IyfWbyxX6wNkh/FFBG+ty75wVnpsxUgTG0aUGaXED1QHksNE7+T0d4njLpJpB/myw26KxyS/v8aOlG+8cq27fukYQXbGzpSHPCea7HCfpZR7FbllvjGlz5gorYoK20YulTQCe3tu1FKfJL5FTBmI5Igc4LiMlDd8EDkuAzRqipftXb1SPNEH8s6IrMolpiCj/MjIr1oqyRJPhN0eOz5WVNveLrt8srsmUWQnSL1L5CdT9h3wfMx6TwXZiogyo9MqZ5rCzj6RebszlnIi2RxfJeJnDI6vcn9xRjtW9BlaiueMl3Ie/bxLAiKilGkGX9WmAYou/my2ucysUktMmatjsX0Cumyk5mckmT0ZPWZeNqWckWxL8ptRofqsbmVedd39kucl6Rg3D2tzArg5vhG7XLbx0iqGlGfUUq6t1ovFYg1fAgfX+4jG+zz+Id/d2zd++pO5Y3Bk/thec5kjBEIgBD5ZAhFknyzftB4CIRACIRACIRACIRACzzMBfl8YDHZ2dlZnZ5ecxzdZlvd7JJX/psneiSAibX15DwWZSyy5adPtBY5yzOs6e80Hv9QdILj2WdJ4erTbXT05QoqddFfJM3Z2tEfesd3umPMB0uyIxPzm/zLHlu3UDpSKJSWPqeiRQu05QoznRoG5fFDx5HM/Hua+UjxZr4QYj722vocJ9ZkCskd51dqvskof2rVcu2fwCDN3x5yw7LSWRCrLiARzp8tdxrrHuJVip0fIMpZdXmGZ6OWzM6LgkHws0SzxtTQfveIQqedc7Ic+prThkI1IK1HGc12REWXKOuesLOujshrzNkfH5/LL/nvwvi2HpCuFmDOEgdFfRsdpoPo5s8q1llO6VNXIMVt03o5LlvVMnshJ56y+sk3bsp+eT0Xh1Xfgd0ErfByPS0Mt51JS5oUvq8T9Q8TgEOG64d3Dk9Pje3dv37n94OFH7ARgD1lf6TeUIwRC4NMhEEH26XBOLyEQAiEQAiEQAiEQAiHwPBLQcGyuXbu2Rjodcv3rKIvfJS/Vy/oWdnZc6UCICBo1Efb0FJUoyhp2f1ywMyWvXJpIOFO3QzTSFaLDjBR76cpJd+WY/F1H+90pUVenRIsdI5aOiMzaZfmiyxiNTKrljEScDRFZRkGNEVKVX6yilRQ0Sq0+cqlJGUfTSzKlWZM3PFQ6IXH8GI2mWFMCVXSYogyRoyFSBCmmnCuhZVVvwNJDI73sy3bst4+gMqpsRsTYPkstT4+OKqrs9OSgu3LplA0GrnUvX7vaXbp8qTs7PSEq7rAklUnvl/N5LW00hb3WakreMaRkCaqJkXC1wcF2d0jGzEgqIkvp1JaDNnG2cjdO5rFip0lFlx8jyxRUbixQ+cSo67hZ6ciFLfmTOpWPDI2IKauccryynlJLSbZczLf3cHTOfKNN6m2FG9xKTnqmjrxb2/ykHcWYIF2mqfkS93w+H1Rut8lkthmOdnl4/6WXrv/VD374/Xv81bJ6S7TGXzFvcoRACITAJ0kgguyTpJu2QyAEQiAEQiAEQiAEQuD5JNDMCWNHALl75RjHcR3Z9F8RvfQ9ooYuz4lU4p4VdqRj32zMVfZYqLQpe2+E0arkWAmyjqWVw3VFjF0720aNIcoUY8dEip0gx/Z2Z90+YswE9sqZJsbcNXKKeGk7MZp8v0kpRRamhYguI8AUNFgY+tueqW+EUy/JaozbpYK2XfJnW0dJ5H0tc0QItXsEmEKKpZUlk7hW7hgt5dnyDKTNmyIV3UbdEmUTE+sTUebySxP5I7wOkGJ7M3KpHbB0lGWYns+OjquMdVbs4ukSzMX8orgplkrE0Zm7XzoG+3B+Lm51bETztWgwyvSRX5AvudaPs6LNWNqqMJOXX27brIC5bb835yEr+Xl2HAoydFm1b79zRSdzLvYwcBy1hJK+e85NVPLGKD7L+v14rj63OcyKm2s7uzUCkuix0Yy7QwTlLQb5p/fv37/x0UcfORbD+jxKkNlWjhAIgRD4pAj4r2yOEAiBEAiBEAiBEAiBEAiBEPhFBNi9kuWN0+n4/PziAAlyuNqsJhVZpBRRuhCypADxmYc5rYxAGrNzosv9sGc+5dqcVpvujAT2L18+6q6eEVlFdNUpyyv3WJZYkVDIswrUQja5xNCop9qJkvbbro3VRUkj5dvS/GaoEwWQ7oQ0XyVjanzINMflrpYe62WLhhoPp7U/YikbxmjU1pAILUWP4oeNFvVSTYJ5gfAyKqskE2VcsrhgYan3lQuMtuuaskabKXG8dwkjk+hmPF9Sfr2z6Q7p7uz4pHtwsehu3f2ou331fnfn9t3uo4ePunt373cPzx91H9y+1d29d7978Oi8kvsvh4uKumIfURZXsmRyzq6fnMdIQb2REWbKssqTxhvnPp7MahmrY5kwfSP4HM8CWBu+B0bMWP3OGFBFp6neEHyMe46ks17LQ2Y02aK+EyPafL5czWmTfGmyqiWteyXHgEILrS/LFXUk2UgPZnsDXFcJOE/rwRjhx3kDK/+CDNeL5T4NXuPv06unp6d/+u6Nn7DMckijTXA6r/7vWHWUHyEQAiHwMRPw/wrJEQIhEAIhEAIhEAIhEAIhEAJPE9C+YDaGm9l01+T4e0iPL/L5NXJHmYeM5ZbmGxuukUpGkFl+eyhplDioDZLxl9hYzrsp9urkYLd74/ql7rVrl7rLiDFzdB0izKbkIxsjUcz9NZ2RuJ/cXsqtCRFYY5YbGkVlxJOyyh0efWdyeJ97XUKGCCiXEyq4Sk4xApp0jFz54eBBlacOw9++841yrEqUNKp6rO6zfa+tQ29V3vxfrb++fLt/Mo4mydpbVBR1/WPy+jEyyjntIpvc6fKEiDKvjSbb252yrHSXxP4sv4TTGbnLRjCTzfziolsRVbYiGm/KHBVbSjE1lJsSMIJiV6KMa5PtOx3HWfLOqddH8WVkmNKpfWWWc2WnJZxDgaFtDBoRaQoyljoiEt1IwPbckdPvYjhC2PF9WZ7uiDjjO6fNWq7qnPnYt7tw2nwx9Tviue3YH/nWNhfn53xtI/PcDRaL+QPmeJfdQu/+9Cc37jFOE/ZXdSpsB8dVjhAIgRD4BAgkguwTgJomQyAEQiAEQiAEQiAEQuA5J9AMBu5kynLHzWCwiwZ5g4ifN8hjtefcSnIQhuSyx6cje8p94DKW8wXRRksix+aophUJ+WfddZZTvn79cneVhPwHLD3cISG9emeH3GLrEiy4kGZramllJarH4BiE1EdrKbtUQyXMtuNwLP2HKCSetoT8jLfMTI2pGuEVR4mkkkG85mzUm0n3rdc+2/lxNzBCy3ObGIKn/QpV4o1nEKhayioPz7bHHgYlg9Zcs4qw3o7ZrXNDVJWybWwyf+TY0eFe95AIsoeXj7vz8/Pu/sMH3aNHV7tz+D0i0uyDm3e6O/c/6j6896j78Y33uw8f3OvWjoFIOILiuiH5xkYs5xyTS025uCDCDLMFcWayXTLpVCtJP6LLpatGlD16uGDZKhsGEGI2xG+an0wWRuEpttCMRL4xN77DxcW6Y4T1nfRJ/4erlhduwHxIIVZRci4R9Ttr/aq2lGeras/ln+iyGrecfEe5wQhhuEDaTQfTwWRn9trFowffOzg4uDGbzX766Hz5sPSYIW/t8AvKEQIhEAKfCIH+H5pPpPE0GgIhEAIhEAIhEAIhEAIh8FwS8PcEbMZgfcySQKTHde5/m8/3EBvX+VTOMaKBBkY1EWlVO1g6U8UHYUoImSXJ4lnah6o5RIS9fuW0++IbL3evXLvcHZNr7AA55BLK2Q4J7+mqllSynBMxUgnqvTf6yKgwo45aNFcTUt57KK2evu6fYXqIvtoKK8pUtJQy6alnjrNJtRbVxMhtcSvCPPvk6TbatS9+pk8LclSuMq5r/txbRlHUi7s+Yss2FWY1Z/OsQdoosV2S+++x8+XRwX53dnJMTjY2K4DTZSLKrl+50l2/eqW7dvWytbv79z6sfqBOH0R6kUC/+mFO9ls7TTKWJXnEHIP5y1w+6dgq+ozzemGUn3OmPDgVXxVZ5mRQfgvuK3qM6yURgG0ejbmCzZxwVvS5u11WrZKbjR0Kk9YRlczRbiyHaCWyrX2fNRbfF8ySZYq0PZap7iNWb7Jr6X98//33brbvpfuZXGTVWX6EQAiEwMdMoP1L9jE3muZCIARCIARCIARCIARCIASeawJanzI/+ovler23M9m5ihi5jJOZokVwKYiZzYoAMsULgT1KMSKXFCEuzVsR/TREnu3tjNjB8az75lfe7L7w+qtEaq0RYMig6V5FFimHmmRp5z3EkEv3anmegUPKFXNdNSfGoIz46uWWQ1RwNUllO2oZDyO4jP6qa3Z35BX3NfImayhQOcOqXcRRlWyTth3XKCqQ+t0Y2xt+tq6qDasYcWX5x2JMbDxjiDxXILWBc4UOUlCpyPhD+8or8/8r11CO5BOjEhFVZFbrTtjZc8kYF3BVSBk19/D8ovvm17/U/eX3f9T9n//+/+p+gj9yxnL/aH7O8kY2Btjb7yZIRj9+L0alKbymU3KIMf/JaId+z5FaTYoNRnx3Zvoi+sujZ+tSyoqNY26Ocw1DvGiV8d7vuGScG03yd4GFthWF5zv/ThiRZn400vAj7Fq9vv0F0WQup2V8gwF1B+vBqr5vUpIRkXdpPBhfZ+fUs7/4y1l3cfGoqlXH+RECIRACnyCBJ/9SfYKdpOkQCIEQCIEQCIEQCIEQCIHnioBWR6W0OmKXRYTHFxBiv4MI+jYKxST9pLlyISGahx8lyxAiiiIjkUq2IFBmSJ+rp4fdl954pfv6F9/srnC9T5SU0UfkmaqP0UfWM3KsoshYeqh4GQ2JLOPMRRMxW9nUCxzrKFVqmP7k3kP95H/94XMlVf1hPNzUp8pXHWpUGcvxUWJt67cy2i7ftRa3JUzRRcnWr+Uej2vbuQKsxk+ZJpIQTcgx85BZrwk0WmOKLkN0fF4r5CoBvnNHcE2m5l8zx5jPN90B+cmuXD7rXn3lJZ4Nu5vvv1vLU6dEahkxZkSf4x/RjnnPHNec5ZqOccoy1wXJ9OWxIILM780xKbv6Q9lo5Ji5ysznpvBy7nOWcvpOean8GlJvxtLKGjSV+10x7c/5GvEnoZpT3Tex6ffjWIbKQI4hfw9onmpUpLRiDxLvAvivHnx0/5379z8kWX9Dtj1vvwlr5wiBEAiBj49ABNnHxzIthUAIhEAIhEAIhEAIhMCLQqBUDRFHJciQGl+ajCa/zeS+QdQYtoLQMW4QHeQga+LDpX7KMXc5NHxrRL6rS6cH3edeudp95YtvdK+//FK3v+vySQWIoog8XE/JMcXLuJLykxyfPGIllRApLrNUqJjrqkkX5QpRU+gUzyWhNDi+tyztUrreKYJM/q+NMleYcsZP1WV5p1FZih3eloKxnzJfvtHsUHBEHz6mOgflbKHoOH8hcMNRgov27MEX1aZlvbZ/i3JtccfQ5mKAleWpzfhVROiq6sz+LQ9gShtpxjioyyxrV8lLp0fd5xGP11myeuf2e90Ht4wm42A+cyLN5uZ/Y/zyMUeZXNyZ0kbcXdTPEjGmHKMbBkK/jpNIMcXchu+vosQcOPfL+ZyxNMlnu0bDTVg6W9+j3MljptizeMm17XgVbCUyqeu7xolhuvSSozHnewAN7Q5YWrlk7nfYfOADkvjf/PGP375HMcPbWKFZI3W0NpUjBEIgBD5WAhFkHyvONBYCIRACIRACIRACIRACLwQB7MWAlY3T1Wx3z8iuLyM2fouZfWFVyxUHCrK2e6XiA7EyR7RsyDtmsn0jkJRhL1067b6GHPsc0U4H+zsk42fnQyoqTMbbZZReK3GUY3W9lWMlVURJ+5UYHwHTpFKTTi7j6w+9SRNKShfciffbl24iUGaJJyW9EES9YFP8WFD59bgGworqTM7ytoIKopx1HadzVVr53DpGVdlMNeRPqpQIKv9jW61O/75KUmdVlShMmzWvrcyqpaHbOm1eSCvFlWOgZZPxtwgzBNV40J1dOuteeeVlku4/6N4lmmw+5zugvIO4QGqVeJSVbdg5impuFBnt2a59tDl59ju0rxXLav0emRjjsm+XeSpAx0SNWcb7HcTbLn8/PIqtrcPPJZQOwP4QXvzkOWOovmhSjiJUkNaSTMPJWG6pION+w/NzEv5/yM6W7//knXfeJTLuYTWiH2wg21S2D3MKgRAIgY+DwJP/Vfk4WksbIRACIRACIRACIRACIRACLwIB9MWg29ndW09YlofS+DKi4zcQHG+6GyESoyUbw4rgNWrJncsqK1cWooz4ru6MHFpffvON7mtf+Hx3/fIpkUbIGJ5PSoooep4srRyRRF554rJK49NcducyQc+j0XappUalhFUTXQoZP8qldvaeSluBRMgYsqb5lFI1vqv6npoOa8KtCS2FnDs9WsTnLj/0mS2YI0wLxk9ET8trJh8PfyrJqm+VkG3biILNGsgkhZpGp55vJZv3vKJZ2qX80r4VR1yXsKqmFFTusEl0nQn9bZsy4neJqtJJIXV0dNR9+Stf6A5Yvvr973+/u3P3TjdHVNoprqsklBFjRoQxrZqXGyj0fRm1pnxTVsmf+DKS+BtJ1kTZiO9sgWyr9zRgveWFOcm6bg8R6iYA9jViTJZxXAwRLvWYMTdRaL0Zf58sgwkrkbeVjqRg4w9rSR/NL4bT8YjUa8s7s8nk7bOz0x/++Mfv3G8t1VcAOXvLEQIhEAIfL4EIso+XZ1oLgRAIgRAIgRAIgRAIgReBAGpjNNjb31+PxjN8x+jrSKLfQmy8vkaacF4pOzhGa0KeFC9GllW0EWZkj6V314ge++ZXv8TSysvdPjtV+ouHkUhGP3nV9zKVAAAgAElEQVS4jHKsANvKsbbcEgnEM9tWTilPSlZhYpRgHtt+69xf+7yP7nKHSM2NIsm+HkdqbZ2KdapetamMUoohpnjfzr63nxoxF7zblrVeBYttx+G9Msuj6m7brvbraRuvsq8fv6VLEDE2p1QSjWclBHnGTKr/2hXTW0WbA+qdkMZrW88xK6OMKlNSvUwk2eUrl7pbN292H965Rz/ILr6bBbnJXCq6RJpNpy5hpV9+KCtrGSXXSzcC2Eqr8p/M1Igxl2X6XKaelY3OZUO7G777XXKGTYkkG7tklffKwFqK6TJOaTH2Eohbt6Wo87tV8C3JjeZ7GKIzncOEwD0k3WK5YT53kZQ/PDw4/MFPfvLO7fncVGQRZELIEQIh8MkQiCD7ZLim1RAIgRAIgRAIgRAIgRB4bgkgZLAyo+74+JgUWYMZ+a/eIjzoN9ETrxhJxbHcrHi1Xo8WSyOLiEDC/Hh2F8nTo93u86+90n3xc690r710FdVGDi2kjonmPZRhRhvVZyvC7LJEikLInFb035ZHUkfpgkChaeRLuzd3mNFOzfaomayvnHFJo95FC1TdbeVZG19NjYgmJZENNglHVBZ1LN/q1QXXjmMb/eVSzRJYzp96jFOpRav1vOUQa+2VlNvWowHK2YZWq4xXG49VOWqJpuOttvVQbemjyyRRUTWFknA8V0663NSIsgW7ViqgnLdjVHbZxUvXr3evv/pqd//+ne7mB+935xcXJa4uKO9wi42c+NiD9ZYk7OfStyU6Wd5Y+ckcg9KrmHCtTCvB6ViQY47V3Gh7s50ScEq38opbjuY481CeWdd25FR9A9xNA9xUgH6Y6mbgrqiTiggsy3mf9n68M5v94P3333uPZP3bb6iarNHWVX6EQAiEwMdEoP0v1MfUWJoJgRAIgRAIgRAIgRAIgRB4EQhgT5Au7GCJiNjsjUeTt8aT6X+DxrhWUWIb9Mh6PUB6YLFaRJRLBV2Stzcbd69ev9Z9+2tf6q5fOu6ODogwQmaZLN9dKj1KUilLtqKmP5cnod9aOogo8Tmlq3zpIgSMAqyWGepQOIxGqva2yqRkjrVo36M/23YJOORYPd++831718Sa4qyvw0VJJVkoq7SA7QltiMi6PnNM9b5JM583uea9146l76eNq1qq575qMsxxNAatjPWM2araoOB1MbGMMlKBRdclp5RnE5etEk12dnbSvYwoU3TdvX23JdiH55rlsc7eXSib6GpCTwm2IlpM4eVGB7bd+igZSg2O7dh852FEF8X5bLq9nd2SXeYtq8FanIvaFKBKP/metIq2rVjz+11WvrIShUyX79fvk79SjOWcqjf5vm8QCXf7xrs3uKfik6MgNbZPHuYqBEIgBP6+BCLI/r7kUi8EQiAEQiAEQiAEQiAEXkQCTTuwsnE8OD09xZ2s9xFk3+D+e0z3Km7M6CEMChFkm83ICKCSZkiWEY9dWvkWcuyLr7/SXUXU7JBI3oTwFeGETFGMaGkUSk12VYdcm8eK60reP7b5dr+VSCVseIReMb0Y75RSiCvebxVSnetaa6S94bAZXdrAHwolH3pGBPHQBuvsqUSdjxQ1vKhn/HDJoGamotfs2/Z57rPHIowb67dnSjG7afO1HQPNPKvCfO4Yaow8dCmkmwK4HNL6bXmplRRYRq7xzhfMqUV08Xw8RSaZ/02Z1ZaJrig0VTzR+Rm7XL7+6ivdjAix+x/e6x5+9FHhnZNLzOHXkkqFGVzMK0fDtKPgoi/aoekmzfh+a9yM137s38OzMtFIMnOUuaOlyzyNGmt50hhwtUW7RBAWUe79BmxPQVdtMRbHS0Sgf5+qbUSbGeQWLMH9iL9ft3d2d259//t/xW6WG3ez9LCJHCEQAiHwsRKIIPtYcaaxEAiBEAiBEAiBEAiBEHiuCTR7ofZBkB0eHnI1OCLy6ptE9vwj/MUV83FxlCB7HEFGRNJmMe8OdqbdF954tfvml7/AzpXXun2kiUnklS0Kp/5okWH6E549frzNO7ZNgl9iiAq1bE+xoo3xHpG2dV9VvykVm+nfa7A4mp8pKVRLNut90zND13tuD6VMqTYjwhRVDokf9Yez8qbGyZOKQLO0ZVhM6vnJZgCtng9b+Xa/dT7NqVHe8dpn9UFZo8BsTdFWgo0yjY/9NTnWSlDKe94rwrRTbhjQ1J3ttvHZAa6JZZjD7uBgt7uCsDTf10cffkhf5Ioj+b79l+wSJNcrc5RV5BgiSw6My2d1LgHnCNq4rauUc5ls1UWUyYodJ5Fk7FLqks2lwo4xIOtM+28kmbtptnnDvsZIjjje1zdCAyUJmQz1pDpgCS8FByYp+3Bvb/fG7ds333348IFRZR7+Hmu5NjBvqhoXOUIgBELg70kgguzvCS7VQiAEQiAEQiAEQiAEQuAFJKB04BgMzA91cHQ8QuCcIU3eQtb8GlLlsvm1WE7Jho8rpMZq1AyFOchW3eWTo+5XvvHl7ktIsssnx5V7zPxjiiWTs3soYnpRomQxPbuRWS1qCieioDHP1mjqOEqgmMPL5YMboqwqYmsb/aXM6WWS17zkw4i2s1AglSGjFYPTfK7M0QtZlJ5KgLnqcuA4W5HSLr6rKv7YPnfcHkodjZe37XqrqWi0pA8vFDaOtc2V+Vuxnvmc8v1clF4enP9/9t6sSdbsOs/bOWfNdYaqM3afHoAG0AQgEJRJUZYomyFHyMP/cTj8Oxz2f/C1w+HwhS9kCzItigBJkBR7QA9nHmuunNPPs3Z+dU43AIoQdKOutRtZ+Q17fHeyGf3Eu9YOVxuXTZvIw0YfNIyxvAyA5Vp5FuGOPHSd6iPMi4rMSp4ozNzeXC/X2It2e0HesvNw8o3P4UzWBVyFi4trvx23hkUuyoS8ZIZb2o9ATMkdr4ZYVqgoZHM/Z+ytdbc2dxi5lgZY6VBz71Uz9hiVHce5xt7xPQeouW/oBSBrL/nLq07fV/T2CrD35f7e/v3Pv/j8xDEpCmBphqt3+TcVSAVSgd9CgeZfLL9FF9k0FUgFUoFUIBVIBVKBVCAVSAW+YQosgBmkpZp1gRk7wJMdIElPsCFImQEpAGUREud9wBBcTetrw7JHWOXWxpCcYzVhv7oEbIJ2NO0r1IJuBM+pMMl6BvM1YCWADe8DmNkWLqKjqoFITT3b2V/Tp/cBYHjmd5SIyfQ5IAigZFvnZKmuMcZdVfXdm5+ow7OLsoJT9Z558W6+Gsd2nvxo8Tq0od+Ynyjtjf/6asawru+b+t5XyFbHtA8/Pquutdfz4/EvrTv6dS0AS0+39Hv/+nb53e9/t3zw7lvl6tZauXF9p6z3md98HO6+GfnEDLl07uoR38x/yjOL83MOzbW6Nus079hkNi5HONQm4USrucWsb71OhxNM+bzZPvRY7U/kQ9NJRl3rNPtRx25vUfc6Q9waDtdu712/scFsFMbJrHYsppV/UoFUIBX4rRVIB9lvLWF2kAqkAqlAKpAKpAKpQCqQCvynp4CUoSKYr8y9Ihxo0fr6VukPBmsAinuAi9+FX3yf6x1rA2EWs+kElgF5EoTgMFrjpMK3b98IB9n1nS0AlDmqDK8U/ryGVYbS0ReOo15ALxP3myes2+5VdxRgRscZjagHHKJuAJsVRKJ1ABvpiPMP2MKVz4VDFr997ydcVT6kjv2KmXxj39ZzjrV27csBQVBUrz2I0uyoAXPxKoZZgaro2d7tmbq0c072Ey4pnkZXUY/r1TrMy4YNDx0qUIpwSeYjTBIEBixarcf+zE9mUT9HAyet1uta+AiXqK+TT/kMb/TZwuT7fK+vbwAut8qrw1fl5OQ0wjTt95TcZOT6KlPykHkf4ZuBn+xH4Det/TNXS5MbzjGt72ycq3u6BiDd2NiM/RyPRlUHJuP7aEslT7S0TOecfso/Jvm3rwHhmXwTSRuLDoVpN+PulHGOkfa01++dPnxw/5RZSCGrEIqRJRVIBVKB/wgK1P8H+B+ho+wiFUgFUoFUIBVIBVKBVCAVSAW+EQpU/AOZAExw+GRLSOanY6idH8CFdS4cZK6a92Vne7tsr22Aiio88ZnwowFEX1dHV5RuNIsQzL6tL1D5KlQhVJLis4BAwVCYwOrbd28+d9zmvrm2TsAdL6AtPqfHuGvqxlzps7n322dRXAf3Os/8frO4jqbUfpkPIYcXbVcvm/5ch86zLon2rbMkxLSut85bHXrdgYvifZ1D09auCISMHj14IPpazdHnju98nKdwMq55Ztq1Wzf3y49/+P1y5+bVMiQ4dr1HMv+dTax7E7P2E4I5BsRNCa8cXcw9co0xWgeAiZOrarAa40293L+DgwNmUHUyJ1msH4bqWrx2rq4tdKSPAJ+skXR38Y65ErZbnYnW49PhfpfPO3y+vb+/f/vq1asIc1Ho6mubcfEqL1KBVCAV+M0UeP1v8t+sXdZOBVKBVCAVSAVSgVQgFUgFUoFvngIr8kNWLuBKfzDcBOLchW18CHj5gOVuuWTC3xadFvgFXqTDyFMQhxCYt0nM/9333i4bawNADSAJWKJ7qYKeFWACjFSIFAAOVqWDqgKdNk4mnVjWb7iHzipDMXVaOWBzeqUnYFYuJECqzqrGFSZC0rVmYQa0FTx5ZZ4xx6NNnKxIPSv5Z8XBIFtc254xeWbCe4dtqsS8HJD/uULnFCDIa+ctmoqxbcE98McOoh7vXbvwzIT74Kz4NtdY7c1QQ7qW21Gvhh+SiD/a+W4F9FjanEMRHEGXVx2Vd8176zMH23UjNxmaM6adC652OHzh1avnnG55HAtTWx1nAjLziYXLb+WAi9xujDDViaaCjBFrYWwGCNdYhZsz2s/K9u5uGTCGhynoRqvalNIjr9ySEy9rwn6AoKdfMjdiKqOOc9Uw1uy3cw2tWCTvxvPF7IB9e3Djxv7DL7+8f1ZzoYUEzgTVfl3xd6BSf0eVX9c0n6cCqcClUqD+f41LteRcbCqQCqQCqUAqkAqkAqlAKpAK/PsUEGzoPsLFY0xcj+/4bwecPAFeBDO1DpADqNIB6GwM1y4cSzWUUc7z2kklBPFTwUd1DdlH06ff4JILqBLOqq+BDdvbxs+bJfoO+FX/E+fNcXQjVbDGrGj/Zqn3dU4+F6QFEZPKxX0dr2nXjK02zbM2MMjiO/OomedsCQCLD/BrTl9zni14NmOOEwx4i1aPutbplfEUZxXPRuMZ7i000FFGG/LUx+pdqrBM1tiM04zvHBxXTXV7eS+wCi1p0Oikm6wLxNxcH5Y7t/fLH/5nPy7vvn2r9MkVB8oqa4NuGQAowVilTbvZpOYkU7tmf5yH1z5r1u5Yjuv4Y3KRPX/+9KK+dZp5NPN0Pj5r5mq7uqbqfvM9dT3N0g3uUneLMQztXZtOZ8NBf23r9u3b/CajnXX8ZEkFUoFU4LdWoP6b/LfuJjtIBVKBVCAVSAVSgVQgFUgFUoFvgAIrKiSMqTRmOZ8OgBhr+rBW8EKA0fJkwqaOkENg03yrg/dGYnJ2YoUpuIl0HwlGZE/mngrIsYI7cUyiBIaiz8tK4Y5aOaFmgKNoCw9h+PAExfcFYKnQrM7xNZRjUH1aF6Ao3geEwVUVwzEZXEwBxaLXCrqcnwq0fUeVOfGFrs81+23R+eW1fQrG/LZRXcUK4sHmJoYL8lz4Z/Is+5jPT8nDRbtwUpGPbSbEM+xSV1V1evXCabbEfVXBIlJEUv0FKbhcuz12mUO9Xq2fupwJGvrGc2HUao6F/F/ui+2+9f498n71GO9Py7/7+PPy9NWrAnzCBUZuMAZybN1eU6Cda3Rezjv2IPQTygHj2FNGpl9CJnl/eHhYRuQfG/Q4qIF2c0SuJ5cyL/LNze2fepaYn5pRiOat39yiRTzkPaXdR9c1UqsNCMXc5Hrv/fe+ffb551++pAGnCNS+uFaQ2ln01Py5eN88yO9UIBVIBX6lAgnIfqUs+TAVSAVSgVQgFUgFUoFUIBW4tAoIGgJe6BrrdbAxFYxGBNYJgIQbfkhAFuCkcRNBMkofANIFlPRwKglLxEi28cOfCPMTp2Cnoq2gBjASr2q/9iF0qonsK4SyTn3uVe3P++bafu1fiONzUZXFa+fZON28jx4BXdbpCOAM+4O8iJTs0jr+E/MF/liC49EiQFj0a4io4Y4qUutOhWnBt3CKcT0n7JTecISR14uTIE/ORuUYaDTGbfUKgHRydopDa17Ozs5wjOnGAibOFsUDC7YIf+z3e2V7c51TQQdld3urDLnf3d0Ohjjs4/IyoRjcR50a/Rmuztu5oEeXtbl+nX1N8cqg0uHQnGALDlW4Vf7oH/2+qy+tTz4vz14ccbplr5wzpyl9CEHVQsTkOH5M6C9km5OrLDSn/0Z/odpkMionx4dl7So/G94NBoPQwBBOSw3HrA60Ct4EqRVi2b+6NSXmz0mc7MsaY1yj2h1cZIebm5un77/3/uknn35Uj9l8s1HTOL9TgVQgFfgNFUhA9hsKltVTgVQgFUgFUoFUIBVIBVKBb7gC4cLp9/u6haQfcIx2S6eTAKkpC51VAU9wRQFlGkgyHpPofa0bTiNhiDm9ohmhfAGpCCkUhISrawV1CAyMbn0f/dCvj5p7QUnN0wVzAdBYmhxj9fp1exvaLnxUwBXoS70HhJHjKkYyeq+2APbFOPQSXI3l2nYFlUCC0TYATizC3oFj/NU1ZX41wyjtbMEXGE1JGKdbTs9H5eDotHx+/0H58uGj8uDxs/Li4LAcHJ+gF1qQvN4iIJtyP+wNQjPnLiDb3d4JSHZ3/3rZJZH+/tUr5dq1rXJ1dxMQSX448ncNeoQ2spYuec4CLpkfzPkD7wIuce161EC3l5qZu6vN+zXzhDH+t94bhpPsys5u+bd/+fPy8MlBWQo4z6a4yLplPCbXGePEaaSxtgpIa340IaNjVp3cO5U5ePm8bG9sBxxDIISpzjvfCwHPz89Dp+pmcy+ZGxvR47exJJ8d9WK7netyYf60zvp8ubzD5N9jXa9o/+DevXvd+w++YH7noWP+SQVSgVTgt1UgAdlvq2C2TwVSgVQgFUgFUoFUIBVIBb6BCujuoXSAF4ZWYsSStGgKqo4h4dcM0CX00IXVvDMEz6oBlVb1fad/q9atuc3gKFHsT08X9jRgiHBK7sY9fcBxYryALNT2+YUj6o32tacKWhzJ8Q2RdMbNXOzPsQRKdCPNirJaVvTtg2jrODievI73q0TyMX9cUhabG4IYlIkcZCa6H01n5WQ0Lc+evyiffPpF+fLBo/LxZ58Byo7L4ekocpCZ7L7f11XFyZGU/mCtkJq+nOIoWxLO6BgCp+cHRxFO+cXn9wFlw3JlZ6PsXb9S/uGPvs/JkxvkDOuXDdxZ/YG6GhLJXHW1KSDrZuOiL+cp8NMxFrrG9Kt7bmODE0dxtr339lu07+As65ef/Js/L09fHpR+d728PDoJF9spkGzRNqyzOtbcW3UxvLLnJlGqu6wbDrGTk+MAV0JWXXbq3rQJDVmj8KsC1Or881ABSF7M0f6o1/K3xIW369zfFY51O63PeTQAtHXv3r3b+uSTj1Y7GTvRXNsmSyqQCqQCv5ECCch+I7myciqQCqQCqUAqkAqkAqlAKvCNVwCyUkPjgESSrj5ggo9WIIpOJP60cUnpHhJydIEbAhOBiDGJLR1l1BaGiE/iG0jSFO/9p0KR1VMaLABDUUugwntdS0Kz6n6qIGaJC0zgwkRiTFs7tuGSOsQEWzGeji5wyWvIhmtrNVTTps6jtjd+Me4D+Jjovob9gQZjvA6wRshmeiyBXs2v1iaMcl7OR+fl/uOn5cnT5+VvP/m0fHn/YXnx4mVNzk83E/KLeXKlkMhTJGfcr62tVZcdkFHnVAfXmOvSYbWYTcro7LxMRuPy7OBleflqVj7/AuiF3j/72c/K7/2D3yk/+vDDcnPvStncXCvLPmn20U7DXxsdG33qeqpzr1mzc7AY2qoLbI1xx4z79tt3ywbhndf2rpc/+9lfRV6y5XKjHDCPdcI6j3HEeTql7f2oga67drvPPgkdZVMqbH41XGQHB6x1vfRI/i9YE/o5L/KIAc1icNbJ/nQ98ZT9ZL/42YROANfYKvokWjR+QwLaHca9zpAm7N/ievvunXvnn37y2Ygd4XFdF++ypAKpQCrwH6RAArL/INmyUSqQCqQCqUAqkAqkAqlAKvDNVwBXEIisNQRODEEZQorIb/V65RXoTAA6FYxMwx1lfi6L4CNgmZCDUEv6AK7UExbNZWV/AqgoKxDlM4tthSMdwFf0A2CJ5zqNBCmretbxvdCmPqv13nxvO+9JgU9Tk+1TRxrTPPcdn4Brs/rc/nRIgZuiXrvTIxRyQY6tGU4xcovR/uj4NMDYg4ePy0ef/qI8fvKsnAG1poAnwWGEefb6pU8Y5vr6Osn6ZxHO6FjdrqndCoBrM8DT2uZGXHvv+x5tjo4PAGWn5YywzPOzkzIGxB08f1b+1b/6STl89qz84e//uNy9e6dsbKyRwd55EgoZObtYJQ6tpoizdJEJ+CyuTQl4xDUauy882MehpqtsZ2cn5vvXH39WWqTCP2PNws+Dk1Py/ON+Q3PDS51nU9yH13tRyvHJYdkd7ZZuf8g4utmEi5OAgr1eh5M7Z+E6w0r3Wnv3kj75+koJCIudjP63YWY3+X7f7QE2dt97770vyUVGnCWBo1jonAPlaz18pbu8SQVSgVTgVyqQgOxXypIPU4FUIBVIBVKBVCAVSAVSgUumQMM6VmhB6MSnw+0AG480J0hRcCp4F44tgITGHU847BNiSG4xc2ABatrkrBKeGHY3BwqBp3ALUTcgGE6vVciidQwPtI3hdHVMQZpV63P8W9UFRh3hh3WdivOo7Z0w9/RZ7+t3vGdc/UcyON1SF/VpEu41nnMcJ+0BRIIV1tzipEcBUpcQxjbfJtk32f58NAtAdnJyFuGS9x8/Ll98+aD8zceflKNTk+3X8EidbIInHWLOrI9DKq4Bg3vrG8YGlmtXdsr1q9fK1atX49NjrOHGehnSRkAljBqT6F+Y+PzpU/Jygbim43IGoHry5HF5+uRRaeFw++jjjwF24/Lee++Utd2d0Ecf1YR3ffQMRx06tldwUvKkw0xV3BfnKW9U0QEuNpZL7rON8jsffhDz2rn+ZzjW/qZ8+fg5DrW6LzrJLAI8c6dNOJVSXQWhfruHOsZ8fnoKUGMeA8JIBXa+F3Z1+K2UAkhE2wnQrLYBGrrnbJYw1blT3xLjCeSY/2Z/0L/H7+oUl9mA/ue3b916+ejh/fMz4OEKjtlA6S+KfazeXTzLi1QgFUgFvq5AArKvK5L3qUAqkAqkAqlAKpAKpAKpwOVVoNII1h/5n/gCXkSIJe6qtsArIFVAC51b/OfEsoKjeAfY8JVAQsjkpwl59L2J2Fs6xwJaCVK8qlDFfpu+W4RJCk2kHJEAHhhTXUjWocXFLOtYbtdF2zdemnfL0zaFX/ZX68VX3Ds/i3OzxO1y2qw9winHkwV5xUi4f3hcXpIX7OmrV+Xps5flF1/eL89eHZRTTqI0Ef5sClQDBvUJg/SEx/X1IZCKUykBXkOA196V3XLt6m65bdL97c2yd+1qJLHXWdYlzJEkYCyCOQIADbNsdTDt0e+1rTVOBe0GHBNCHbzzFqGXZ+Up4Ex32QIw9+rVYdmgn83+emjquupeyfwquAr96a8Jh617JLT0PV+NppDFAS6027f2yj/9wz+ogOuvPuawgSdl1AM0YSYUkrneJbpxHii6oRlwy71eub14tgwX2fb2NnszLwO00EHnuO6FWp0CtQR56uWhAxFmydzdS+s4Z75pcvEb2QCqvcv9jM8xn895e/327bujj8NFFnGWX4Fj7qv9ZUkFUoFU4N+nQAKyf59C+T4VSAVSgVQgFUgFUoFUIBW4DAoIZ6JUaCRUAIAYt9YDRPDfDfh6ACANTCrADj1FFS3VsD1dQ8KZmrSfAENcSYbV2c5QScsCoEZ/AS0CaukqA5LpY9JZ5ImYpNKKfjyxMiAb9WeAKqFJdZDBUujTd5V7CXmqwwwcsuq/riP+AoE8R8B5LVdOJs7mrPV0LAHuzDkm6FlMySvGHM2BNh5NSJZ/WJ6/BIo9f1mevCD5/mefV8cY8zTh/gSnl+DHUyh75OrydMg7t2+V7fW1cg1X1z4gbB+n2K29q7wjsf4aIZfAsB7Osg5OO+c0xy01OwWw0Ue/MwioN+iuxQmbXfoROu3sbIV+V6/tkgB/XG7evFnOT0/KfEKIInM1P5jOK8GTwKk5jKCBZcgTeun6U3/+RNhlC4joPiz45iLcZCwN0Nct13e3yh//0T+Jvo9wr7nOs/ExaxiWUQuNRjjsGB/56K660gzxjN8ID0fAw9OTI+Z0FejHKZ24DWex//DAISdWnnOip3nIGDcAGapHDjYnwLMunQk3ec/0iJ9stQZc7iHEc3+NbOFgMZ/d2d/fb/3is8++5Ld1Un978YNSryRj8avJP6lAKvD3USAB2d9HpayTCqQCqUAqkAqkAqlAKpAKXCIFhBRCjo6Z6UnQD5joyU4EGRahCyCm1QAxgctCAkMxPNAcU3Aj6ASNYGsiMAGM7Tsr6CXsKitoZsoyYAghmiaaxz0lwAFcWd975xLP6N9njbvIZ9437+J+VceQvABqwDHwDTOpKK9pY3ifkE2XGT6zGMPQxDGhjCOgz2jlGvvs/qPyAkD26Omz8srTKMk7Nmfqc+rOAFv2sUGI5CYOrqu72+TxInQS19Tdm7c4eXI7EunrILMOeKgM+jrEhFiEJtI+cm4x1zU07/SEcqdlABSbngOscFV1yWHWQU+qxFpd74DTKwVhW4RlngGhLvK8qTjv3R/XGTKis/fgpPgWEHof+htuGRrW8FCE4h1z4p+6d0tOy+yU3/nut8sDTuQ8Pj4um4SBnk/nuOLsj3WMRYl1T2r76jLsdfoRZqmOG2i6QAMh2oJwUWXhB2gAACAASURBVLfecV2DvyHn4rcHGLjXPp+xP28W5kz0a4d6U36V3Q3ekY9seYPnffZg+e677z7++JOPeeyalv5W3fgEZG+KmNepQCrwdyqQgOzvlCdfpgKpQCqQCqQCqUAqkAqkApdFgfBaBU0SUIAZWPiS2L/lgDDFPh4euMMqHM+XHEVorjFzSAlcBBzVhQUuIdE9cC3u29rBLHRvnjAdQSaMJ9YyHgtHAmRJc/gYStlmfAGKcE141RvgNgKsWEAxQJbgZ3HvLBdAFfsVVkGI4rl9ykgqnANkcT/nMAF5mVDMd+bhWhK+6fynPJ/gXDrFnWXy/c+/fFAePXlaviABv/e6tqaczigOGo8r1BkCqrZwhG2RJP8dXGNXAGS39vfKdVxj64RNbhBmOegyL9xWLcboA7uwsEWyfcdUZ+fRBY650in5xIYDINHUvF6EogKrppBG86LpwIu1Mr4naJpjDTtd5DcT9mFDi7507NXQ1woEna970GhMWrlYryKFo85OeaaowZToR5eeifuhTDj3SKYP5Hobx9rLtw/KGYn7nfd5uAXZQ/br7HwcbUNv+nNty647V8hDdhJJ/wVfAV0BpNZzD8xN5txj/tRtTvLUMedvYU4//g4CZHIt/Jo5z3nZ6HW693g35/OA8Z7jImsfHh4CWWfl6OioNQPKZUkFUoFU4DdRIAHZb6JW1k0FUoFUIBVIBVKBVCAVSAW+4QoIJDxJsdsjT1SbRFjt1iZgY53nRlR6eiHRiW14j5CjQinDFYUiFsMqzSHmrSGSU+GVoENUZZ4pkRdj+AToBjyyFcBsBYrAcNFvFweS+cZ0PjmOgEfA0uLYAO8hKHGv/yt60A2mS4x3dV4VzMXYPuOd40pXYnz6sl44wYA1U1xRJ2fn5eGjxySlf1we4Bx7iWPsmETzE+GOPZhri/mst3q4nXSNDcv+7pVyg7DHu7duEFK5GTBoCweY44AISaZPmzbuKWxnI6CNYEuYKGQa0afz0zFmWcMRNh8zDnUMv5zNFKdN8v52mXJQQOQqM5QUSBQQjLfCrC7zWXj6JsCvHSGaqEKY5XJRw1vDJeceuH57REuLe0Ql/ugWjO3lGXN2b3jWZXOG7OH62gAH3KDsctLmdcJGX+iimwPwhrj+znF+wf3GQD37VVNDVYVe3gu7RuQa0/XW4TAHD2vw5FLH89lo1I26sRfuSfxGKmSzvR/23Zm37Ms2wMpNfpvv0qbX7fRa09nkF+i5/Ud/9Ecvnr14Wn7yk5/EWu0zSyqQCqQCf18FEpD9fZXKeqlAKpAKpAKpQCqQCqQCqcAlUADw0jJxPHDBMLVBt9VZb3fag9FkFGFrOLHgLfNWPRUy0FZ1+IBUdGDpRmoBOZY4eSbCEMjGLACVFzX/WCdATQVbsjHD6UAmpcMjgYhhmsIoAUeFJAhv3xTdabK6yCHGoxYQRyeUoXvBv2gjCBKmWVq884V9GYrIRbwz3M/6gpyz0/Py6vikPCWU8gmhlEcnJxrkIlfYztZWnMY4aU1JXo+TC7DTB15d39nhNMqtcvPalbJ3ndMot7eYdxfgh0OM3FriugmQyiMJjplLAxAD8jGwgMzcXbY5PTuM+5NDQipxkK0DotqTHoCxx/sh4ZYcBABUmmtzQ98lkGyGG851qq9rM/fXUpeZrBEopylMAKmzLHRAaOcyA4gFKJPUAdd8H0499Pa5eeCiX/pU0+GgW65sbeJUI8ca+7pFiKWdP31xiA6eXKq81ZVmiKwwzj6c05yXOtoEW+fn52W47pwApYR2Nm6x9cF6eXn6Ei1wy7XGOO/IwRYzXkEy1sFesM1G+y6W6s9vglxky2tUG+Eoe9Rqd3YJvbz96aefnvzZT//0FRMyZnTVS3QXN826mhf5nQqkAqnAmwokIHtTjbxOBVKBVCAVSAVSgVQgFUgFLrkCQATYQ4CpLk6inkwCSRpmQd7+lSNMAkOp4MccZK0y4WTDBc892XACmJoAQkY4n0zuHmFz1J+OxgGoAhAB0PwWggE54roHMBoQiuhzc6H1CQ8UZuEYgpEZKmm4oeBl5V6b6EiqYM1pOvdmXh0hkBDJvFpcBpzCceZ4OqWcu/Myqf1kMgrXlYBpQLL9ifOYsGzq9XGtdQmlFLatD9fKVXKL7RFOuXdlO06m3MT51RUu0bcAb0G9MVDLfsesv4FjjuU6BDWGPgoChXtrONF6uKvi9ErenAG4+oQfrm1uARlPS8f8ZbjEDBs0kX8HTcIwxl7oIHM9hqDG2l0+zwIG4mFDqcLBmpAp1v8aGq00UIvq6hNqsVili3cBGIF9ZS7M6wQE3AHchfePvjyMQBon0Ds+AeDx5pQ1B9xkXrYXlk3Zn1NceBuc5un8zClnUQth1xrAzZx1hrC65wLLgGC8U7fVbxFzXJxoye2yhU6d8flok3o9/jdhLzkMs/sOqclmd+7e/ZsH9+8fxiAsZfVtgv+qz+pBfqUCqUAq8HUFEpB9XZG8TwVSgVQgFUgFUoFUIBVIBS6pAkIEoIMhlPqN2gAKLqQkspUIB6QK2MwPdQKixEtBRquc4MQ6n5BEHrhk+OArnFTPXxyUF5z+OCOs0JBLk8pXeAKEA6oIRgRbA8DJNsntt7Y3CdnrlV1ObVzju4NzagBAGeDaEqBwNmI4oYREghRdTRElyHwEPM5dKNbl2zBQx9B9tuJGXNbcVlqvnLPkTLeYcx70WmWD0xXxWZXJOVqQW+yYKmsAqiWQz9MbDTH0s7u9QcL6IQAPp5faCMOAfwKh6WxM+wn9z4E/nlZZDxpAgLh2nj3gktBH6Hfw8oC5c7Ij9QwhFCat4eKbAu3WN7boh3xlfdYGRBP26STrMK6hrEsgoO+bfWEmXAsvdcjhtgLuCS+ZStXGCwtrt40SuMMVGvI49tl7AOXKGeYBCrvb6+Xu3f3y8ZdflhNyjvXYlxZQbZf9ch/mUEodYyP2U2ecCfcn5FSzP91jAkGvHUdganin4/dxqBnS++rVqzKi3mCVzF9HnCdx+tvw94KLkUt6mLcW5GPrund+gKcjKnHWQesG3+e3bt36/Omzx4czDlqgtj8KO4mx/c6SCqQCqcCvUyAB2a9TJp+nAqlAKpAKpAKpQCqQCqQCl0wBAQagQaggECOaknjLdrsPKOsJM/g0sKFlYvwAFwAPoYcgCj+TMW9l0R2W8/G8PHz2qvz8L/864MTB4ctwDY1J+u44ESLIQJFwP9qT6wooNCCvladBXt3dxa3VLzubawGmhGbmw1rjWR8oNuBe59ECOCOgWfKuQh55Xi3V7SQcAxrxyDWYrN/iKZdxT9twqwFkhHBCshnOse2NYcx3YziI+us4pba31sjDtRknUpqE33Zq4OEF5ySj98TGkbm4CAcUMG2sb5cNXGAkjceLB+BjrB5gyzxmSjnHLTX1hEdBD8ra1/HhEaIsAiptEt7pHAfce+iBJGuxHOMoG4ZjrMX6BUg6regh5ml99W0Dt4SYEXrqO6rO6L8L2LK+hxrE/AFuHlTALWXlQuMq+rA9186VZF/syU7sx5OnL4Fn7DdgboETbJcQzHpAg7U5sIF8bq7FObtGc66dn57FfacjOPS3VF18NA8geHp8RrtROMgGHMrgHKPUia0ul/G7c78DykVuvOVN1nHGgQsHwMbHQMb+lStXytPHT2zjqmJl0UH+SQVSgVTg71AgAdnfIU6+SgVSgVQgFUgFUoFUIBVIBS6ZApiSwn4EV1nAm9q99nJh5qg1OQV5xyKrPnyD6yksJqBZQBzzXR0eHJfz6aycjWfl/qOn5S/++m/LZ19+Xs5P6imQ5tFqIJb8w5xYryFTu7w4fBXvP/2c3FcmwcfBdR1YZg4sHVs7ALRNgFUkjce9tUlye91HEZoIabMvrVLCk/rNRAExYT5irkIXTUXOwcMAmHjkw7K9YYTr9N1abjHedhkBdebAI9dIrGnk21qj/wHQR9eafU05zVK3mGGB56NJGRMaGXBIVNieldPJohycz8oWoIsYwJir/e2wnh5hnMKq0fgct9lZecaJmXNgmSGKUzTss4ZjwJpwafvK1ZiHYGwNd5mhli0StsEuI0+ZOd9eFzaKzXKcJQ61lgcEEGNpSKnQLNaEIAJNT4RsuZmr0gLq6Z57/YQX9NUDoPVps0mY6d396+XF85fl/hNSffVqfrTB+gbQEE020Q/+eMx+O2/nEO45tDo/xw3HXvk81uiBAsJKc6DhRNM1NzkYhaNQQNbjkAYdhxW0AUJXKeWwiulsjLa8u0Ko5g+Z5fp0OvlZp0tg6XK5vnft+hqATGeZrVbLqWBUgJclFUgFUoFfpcCb/yb9Ve/zWSqQCqQCqUAqkAqkAqlAKpAKXAIFhBkWIBMnVBKUR3IrQFOXax1kfR1FPKx/uG7ARRsiEm1p7kmG5hx78uJl+fOf/1X55NNPgSlPw4klRBJgCa9kMiZdHxGO2O1No68eObamy9cnH55y8qFhd8+fPy87gDIh2eb6oNze2wMw4eQCYjkH+1onh5fJ7IUfurTM/QXbw3ClA4pQO9bmHP0AWC4sRQIa5yRwibBGANRkY3IBdwy9dN2GV5rNyzxmAZ94phvLa0NGdcWdEnY44b4/BGABCzHQlTNCBk8evSDp/1lANHNxCQUBOeXOrZvlex9+UL7/3e+Q32u/3Lz7Tjk7OijPHz8iZ9dxdeR50AFA6YwDBGhVNgFGY/okwnAFl7BfAb3YFL4aAFTDJZdmz9cZxjuvhVCGZxaAmfBQx1rsBYAqtHGdPIvwTMMwWUMLgCcMnAD+eoy5TqjpO2/dLE+fPyuHR2flhJBSgiVLi3DUzQ1DLcFrOAjn5lajX06XZH9r0n/DLQ177K5X1x0TCd0NzfRAB0MyB/211y4y4JulE04zHHQ1d1tL5x/7vjAUlX0bzGbzu3y3uH+MVtdxC761u7s729/ff/D06dNzd4xP/XHXa7vNkgqkAqnALymQgOyXJMkHqUAqkAqkAqlAKpAKpAKpwOVTIPJxsWxAE6SEIEHiAOezGfwrwAvOnEXHXFdtoFNAI2gKLrOgD6rlsxNOf3zMKZCvAGT/7q/+ujx59hTAMwLm0C/gyhMnwx0ENDk9m4BWSOQPXBJSTRbc2x/9mN9KwGJD81qdnBFW6DUnLVrn6GQ92gnkWj06Bw4Je1pAtzkATFZkPaiW6ChgU7AR+paWWCQmzkdwZC4vP4YL9oBA20CZgG8ApRkuMfOLuQYT3xtaGlBsPGINfABjx7ijTllHi2MaH+Oi+/TLx+Xjz74oLw9OgEScZnkRcgiwYl0muO/9xSel/X/+y/LW7evle++/V/7xj39U3n/nrXLz7XfK6fFRefzwQVngJHMd5vDiHEfykBFmuqH7i9VwqqYAr4frqw08cn0CP2VjmQG9eOgi0RkrlVAslHDPqMc/ai0ujLBTSSP3AQFJIiZYDPDJVR8wB5laOfq2yrfu3SlPn7wM6HeC+802XSDmJq6/yTpzZt5zPvxSYg/DtcX4uLxKbw6gY84xUefFOsi+xj60ywBXoI68EW68Yb/mrKv7yiyZm3sSgNN5s88VbsYBEFv8Xt+m7ivAZYd6k3fvvfMS0Hh+Sl68aOTvQZGypAKpQCrwaxTw36RZUoFUIBVIBVKBVCAVSAVSgVTgkipQIYiLD5NNe2N9q0MIHDxiOeTdtyERv8fLdwEPpkiH10hPlm3D8yw6yAQsgqgFEGWdsMePP/qoPHnyhKT1Zz4lFxehgTh+BiahJ29WQDOeD7k3t5g+ryFJ8g059L2nVJqgXdAlDhLMQXiAJ5xwuHKACY5MrC9AaUc7HFJAH5Pz87/os84KqGX4JfMMKCZ84x+hkq4k1gdoqoCtzxzbOKY6DBx1+eNJmOY8W+Aim5kzDGA24XN8fAwQPC8vDo7KGTCos7ZdnhJa+L/9X/9P+ej+ozJpDcqL03E5BKCNNGT11kheT24tPh1Obnx2cFCW9DvGVfUcoPj//es/KR998kl5+fIV4Ze9ssOBBZ70yELCJWd4ZEfnWMyvArHYO9bT/INokVvM53U3+faaj6U691ibt96wNoGT73VmCdgEgLaOOqzZC7W2Ttf6wZhahFEeEwJ6HOxrwhp66s60BJo6+IRtDjHFOebvo/I3YBungJqDrUK9mFboTfUoE+AY+cTYW/eCesA5x7eDWAcVnSe/RR2OsbeCM6Y35H5ICCnVly+Gg8Gj4WB49AwHYl1sdJ+ArMqcf1OBVOBXKJCA7FeIko9SgVQgFUgFUoFUIBVIBVKBy6dAAIj25uaWUSYYqjrrQIjvACX+gPt7JnvnQ3BbJGCXaQVgEn4Y7iY8MpeXSdkfPX6Ia2oSgGt7a52QSHJwAW+2gGfXyCl2++b1cu+tu+VdnEjffvdu+fC73yo3ruyW2+S3urK7Wa5f2YlE/Vc4IdETJAVsbdxegivdU8IbYRsTApZwEiJAyUT5ghfz1rdwK+mbCsgG0OFxXLunusZgZQFoTBRvSKHuMRPKG4qpp0oQUyEZoZSEOAr6poQTLgBBx4Cto6NDTp48Ks84ffIcXrh57UZ5eToqP/v4F+X3/uiPyz/55/9NuXrzVvm9P/jPyzvf+g4nNW6UR/fvRzL8KSGI27tXyv/8P/0v5YyQywnus+tXr5Z779yTKRFS+iIA4+HhwQrK4Uxjvmu4qwRGPcIXWcXFP+oiGDMU0ef+L3xysYaaw8v1RK4xn1FBkCgYAy2Gluwz98A3V88cApQJQIVm1Fc/CBr3JusHapIjTDeYp06eAgU7wCuhVj1RFOcYdYWZhtXGoujU6NwpOdG6nD4qiOyYXwyH3sJ3tFd/1+BcR4TXdjnUgHz7sXadYv6uPNF0pkWOSizTeUrOdDd2+WVu8Jvt8Ps85O2XuOUeXL167YC0ecvDw6NQxVXwyZIKpAKpwK9UIEMsf6Us+TAVSAVSgVQgFUgFUoFUIBW4fArAFwJQAB66QJMNPtvYcTYqjpB1CDqEGdarIW8BV4Bk5qgymf2LF88iJHANaHXzxl65ur1FaN6g3AUYXQGCXd+7WsgRFTBNJ5n5sEZxwmEPZ9kkQhY9DdKwQnN2aR7y+wyQtATaOP4AuCJwE4iZV2vECZKbkLH5gA/crCvsEZTpgAK0VGikS0w/m04pk9HXdeiJgtZU59UKFBnKOcP5NKW9kEd3lSDr/Ow0nGO6vI5wh7X76+Xq9b1yADj7i48+Lf/sv/oX5Q//+F+Un3I4wRd/+hcArhflys5O+a//2/8uQk+fPHgIIOqXx48elwPcV//9//A/ls8/+uvy+IvPytGLJxwAwG9uPimHL5+V9nwcbTZIjI+KZYjrbJ1E9oYvLgkL1VXVZr66pzpwohl5vDhzNMJN1ciPdfyOPRIE8s+CPG+G01oVdhQ/crbywpmnWNWRRQX7oN8lhw0IzQRovC7rQLp7t26UU9xz5+RHe/7qlPxxOPUAiUOcXws6N2m/4x7OT9likZ2LY6/Q0HxvXTbIuVEJUEa4J+v2d+W+WUbnkwCvHUJoddI5fqzVvfJHQTueLYWyALLWZDxusVdbgLV16q9Td2s8Hm+8c++9s2fPni34DTF52mVJBVKBVODXKLD618+veZuPU4FUIBVIBVKBVCAVSAVSgVTgG65AOI8gFbiyBoPW+nBdbNEDXlzj8wMSb/0YALE3F4AY67iArhDeppspQAXtAqjwPlxdVNFB9MG33y/f+eD98ns//LD88Psflu9+C5fY/tWyf3W3bG0My5IcXm1AlPnGNsnJNQRweS1YGQCyBriJvG8DwPrc7+O62iZJ/xr1BsAST5wcAk/WqO/3EBDWtR2QRfjTo70uKYGOIZRx0iP0xdC+cE/5DWgSjnWAVj5nVVaO+p4oOePAgRkQ74zTJEdAOkGdn3NyipmMv7+5UY44sfMzTuz8x//FPy9/8E//uDx49Kw8fPS8fPDhD8oXXzzAcXYM7BkRMjgsB7jChFFO69OP/h3rAtngtLoBSLxzax/XHSGbTwjP5GTLHfq+DYTqMr8+Tqqdne3IubW2xqGiro11Nt81VJS5x1by2H/YJv+xniCKJhSAmS4xxg+3mM/Zt3jvxCgm5ud1uNesC4kK55ZuPT+85pHhsdVxNgUOTibk+eKZJ5n6WzDM1WozAOMpzrsAq3VkYBeJ+gmN7XUHdk2X5p1jPuyd8/KP4O4c2Cb8Mv+Z+2XmNOe2iBDOes282bKYeHsM0KTthENYnzGVhzjanjHuUW/QG9Pf7OXLl3bu5PlkSQVSgVTglxVIQPbLmuSTVCAVSAVSgVQgFUgFUoFU4NIoYJghRXIAhNlprQ3X4El4kVqtHQDDdwAQP+B6n9hK4ceCnGPcttrmGxOQCUQEIEKMoQnu19fLB++/W370gw/Lt9+/V+7c2C9XtjeAZ56CSAimSdg5pXEGIOuRa0xn1nzGB8AxAYqck9tqgoPs6PCVhAUgMic0cx2QwwmVgJcNnVSEG3qi4nDYw80ERAGkrNG/37rKBC2RF42LAEQr8OXpj/IRwyrN6eW7doeQRcL+ugCbDu0jNxbrWTKuLrIxjqc5UOeUeZ3hdNPJtsaJjV1yaZ2OpuXhs5flh//wD8ofElp5jOtpc2OL0zzn5ad//vNy//6D8ujL++Wnf/Zvw2E3wRU352RHId46kMgTKwVwf/WXP4VDkseM0Mc1qNlbt2+WvWu7ZXtzs9y4fr1cu3Y1wkhN7h+kiy3rckpnm3m3AHsRKioI4x+dVj4L6MS1OCj2h3f6uNi4cItV+AWYUixKoCMbUdxbtV7CngRiOuhaurx4756rrTndrHOCe09IZtJ93/HbiLH9XSi2/a5+Y9FPuMXol/xg9A3oW83VcaMt3/aD+4t1AF1xq+ksEwI6L3ORGY5pSCfP4XsLtpHgTCaKc2xBOKZZ/0+o+IKqz+nrZHdnZ/rw4UP7dTVO6aI4ZpZUIBVIBVQgAVn+DlKBVCAVSAVSgVQgFUgFUoFLrYBQBIQB7Liye007jgSM28hB9i4M43cAC7cMk5vP5iAKzk/kdMuALrSpIATHFhBjF5fTvdu3cIu9X955+2a5ef0qDi/gBmCFEzEBXwAiQhanQKYFOayETj4fC8ReHZD0/YjPSeTmEnYJcQQojBunVnJLKCGYB4ASFKa1iHGdu+MLUjjNkI85yXQkAXl4xwueAVq4Foj4XPdYfBinAyTrmttr9c6fgydaLuPkRYEezjFO6BTK9Mmj1sUNZj6tUxLK7929V374e79fDqmztr7JSYxr5cbN22V/f6988rcflfOjA8IlZ+Xk4BX/8QUwYt0ToNsmoZPj0Un5Bx9+h9xmZ4SMlnDX/f7v/rBc29kMALjJWFs4ydYBYzU5v6GjQD3WCAqLb59X51hdly4r3qzAGdeuifWIygKhiYgEYIanCsS4DkjkznofpeprPffA9jrN7IudRAeuA0R6eAEwi/1z1CmOOyFc9AMgs13tEccd83SfPNzBPGLmMeuzJ/zS4jfkWLW262gB3TwMYRRgUCeZv4PanyCsnrDJOLBOF8gRq0QF00GPAxk8XGKOLi/p8iHzej4YDMf93qD14sVzVI4ZNQulSZZUIBVIBaoCCcjyl5AKpAKpQCqQCqQCqUAqkApcegWWrU6739ra2oJhBESChyx3AA0fABh+MJtPbxvaBijjgEDSqhNiGRAE3YQZcQ1A2QQO3bm5V95961a5Rdig4Y9tYIhgytMMTXYvbDKEMJxjOK2OD4/KK0IPz07PyTsGaAFcdQkp1Nk1BkKNgS5Hx6fUOeHEyENCHGlLHq4xoInJEHoH7MFJpatI6EOInZwrQJLwxU9AJQCLRYgWrivzkOEoEzDFtwAm1g6QA+548qVERseXDinvhV9MEMhDwnnmsLG1U771ve+TE4zw0OF6vD82aT0T2NrcAn59t7x69rgcvXxeRsDAfguHGPGfV7fWcKYdlbdv467bGpbvf+fbQMV75Xvffg8CyFjk4yJqlHxeQD36QvW6Htfn/J1zrIN7YKALdk1ei8NchzrolcKEBVyiCt/mjTNnm99sWugR0MlrYZjCoaf7JUeK24Bk4i9DHwVm8fswdVzU9wTLmbCTPZq4x5zwOQZskRyfCgUIZjhlzRumy8u8bkJRgWaPZP38PFa6MyQDOhXnYd4xfw+28YACc5bZn92qgbnhOmhpXe6lcq7H3+WAZ300G3H9mOcP+D4xf9uzZ097M35TsVhrZ0kFUoFU4A0FEpC9IUZepgKpQCqQCqQCqUAqkAqkApdOAZkIjKHfG3YIsRQ4zABEJum/AXj4AW9/CLm4sXKKYRgCpnnEI42oA2vAFTTH0cO1R1ve3L9Wvved9wE/m6UDzQgo4kmQ5u4iHG98dl7G52fl8PCwHL46Itn9Od3jIgKEDIEY9B4hik+eH5SXB6flybNX5YA2E/LtTwBXhwCoA9xc54CYEUBmAigx11WHxPyG4Qn4InRPUEZeKx7Gs3pSpa4xoJhgjPcBxwRjwiZAi7mvZpAfYZCgSOTiaYvCJ9EQzjmeVEAkLNvZvVbmUKjzsxH1DPlcAwwCvTipc412c5xiP/7Bd8s7t/ZwkD0vG71WuXdnjwT3e+V3v//d8sPvfat8e3WSp0nvZ2NCOI8PI4fbgBDSCrJMkM98VNy50i8XQEEgGc9dgw44LmINAYx8rkuO7yYfmHtlN/U/AOmT9bBiu+U51y6WOtXJ5TXD0Ec854YqoYfVbBkuPquxJ+c4yEa46cbs8xHzH/FNV0yJwxTIGSe47AExl05ASEd7e+ms9kEwxmTj9xROMefD/owAbVMA5RCQZi4298K2M0DdGHgWjj6gIPvOdAyf9GcYoM/D6Oa4Hp8R0vkLrp/pQjs/P+scHx8zMyqtinplSQVSgVRABfwXR5ZUIBVIBVKBVCAVSAVSgVQgFbhECggFAm69XnNALyDDPNxKUAreb/J6h8+a9QUynjKpjA4TWAAAIABJREFUe8c6TXtPfLTMcIPp6jk7OwOawB+AY12A0NSQQhxjU4BWi2eeTincOMQ5phOrZS4q3Fxr5BnTMXbA8wcPn5SHT56X45MzPvXUwzY5xoQfMT8oj7nHNkjaf/P6ToCtNZLmDwZTksf3y7SHC0rnGq63FgBHuGeYp3MWewnzFpIhKY58RMAHDPJ9aAPEMSQz1jYltxlz67GuAYBsOj3iA0QDvh3haDt7/qqQdr6UB49LZ22D/GTrAKKqiadzHh+9wh13XLb7y7J35zpAalFu39zHPYbL7uYNco3tRLjh+ckh81rguuvjrtL1xtSY5BRgJ1hyXo4p0hICSrsEe/wpoqGAXF+DPcItcZShosGEqOeplII3c7u5Xh1qfvuxX41zXkMqo57jSpPYqngvWlJFi3thaKpg9fHjp9xz2iT1zCc3A5wiYUC5NvUGwjD755r/lRF7rYuw0yWvmvNY/a5ir7h2jkKt07NjTjY9I/fcRoxpPQGZ7+KETeZJ6jFMc3XxWCEJj53D3nrbhNneQC3h7uf8Ns/2rt9YPnr0SA4aJfa6uamP8m8qkApcYgUSkF3izc+lpwKpQCqQCqQCqUAqkApcTgUCgDRLX8ECgYPAwALEIMquzTGDpU9d3WQVmsRbr1egKoCH4YjVkST4EIAZHtcD5phvbE4o4hIYMgOuHR/jGCPPmHXMUDWjfUcH2rJTnr48LI+fvyx//befkc/rHDBmmB78B9fQs+fAI8iLoZRCFhPGG765O1ljLhCd+S6wbB2XUYcwz2EZMBFhnvWrg4z5TWJEeJJkDGAGlGt0sE+vhYA6lhAioBvRpIwH2GGuPRxMJ+Zh0zGFs+n06BwANCgtwN05J1meMt/RDG2oKyQT4lgEQ1fIN3b7B9/BzdUq29ubZY/cbLdv3CR00JMc0Q99as40whGZn3m+XPyUUMuAOPTT7I2AyPl95Z75W+ruxSXv3ViBn2urcMvTRc3JpmauVyCn789if+5jU2r/r/fdPgybJB9+rHG6qqvjqw8k4wTUAKPugfBtBBTtCSbZlz4axS+EOe1wL2zzxE7B6RqhqK0WYaLC0sjSxsEPzop5dokz9bd0Cmic79AX/bieHmMu3aspjj8Ardpt9NdZEl40pJuwS1xr7hug1D5r2ScU9NHa2tqI9SlMFDXIkgqkAqlAo0ACskaJ/E4FUoFUIBVIBVKBVCAVSAUurwLQCYw1AAM/AAUdZEIKIuigHBSBCfcYsnQgxXXAIq/NDyVq0UF2QvijRZAyC2AE2ACa2E0FaOSpwoE1N8TRsDeg04uHj8qnXzwoB4CxznCHcdaBSBvliL5evnxZ8COVHnAFjkQy+5Wbjf7OgW9nnBx5ghPpnBC/BZ43Qy8FXRuArXB64SZzbD+Qvupu054VM3ZOq/XwX0arpcb6XIOwZzYCVAn6AFZCm3US8QvNru4AmoA1hhNy+CcZ9oVr1VtlEn1dXX1OqlzHIdcnIf2ALPzDYR+AR66yCBk0TJGQTSAV3eC8ElShonPkH3OfRRgjOnlipOhKrYVbbU6wjJxchluuiho7v5pH7TUqW+0n49S9jd5dC+2+jofs3zDVmIN0klLHjMvVdYWjahxuMF71PFF0APhig0eEWwpEXY9gUUDq3KgeukEOywbrd79OgJbWHzgbHWuES7qGKXvF+ZSrdt1wHPq72gGQeQiDc/JjcUzhrnsU66/v+J3OhbzbfN+k2h6fl6zr/Nq1a63nz582y39NBO0sSyqQClxqBRKQXertz8WnAqlAKpAKpAKpQCqQClx2BcQMghLhgniGSx+Z7LyBZFOuBWgtQg6NTlzBiVVIHoxHSOFzT3Y8PKgOMR9o4DJW8Gw25oK8UWNOhCSZ2AFhk63uoIyXk/Il4ZQPnr0o199+t/zox98j5HItQNjJGcnxcQ8dPH9Wvvzi03L4/CnwZkHer10cSS2S3z+N/paba7iRgGVAMnOSjcbkq+pOYj0Y00pvarJ6JkK4nwDMZP4t5usHbhPFtftO6ELOqgqIWE+bvGaLJr8adQacXtkHTvltjixC+8ounXiwAHyH+dInoZ+uVQhmfxu6xLgX4sjlhEa6u9RLWS0Kbl1vdUzpIPMZD/0bxdBFKwjLmpxpAcOYlzm8XIMfQy6bvrx3DL9rf3YRvHPVK0/RIYqD87HeUotXFN5xUigzjnxnutqiNpAyFsxz4Zdr3WVfvD4l15y/BxrWtTg+UGsA3IKZol0X3InLDlh4Ph2Rk47fAsCRt7SvgC6cf/QhhOvzOzk/P8V9eMwhCEMApTnXBGkVvLkex5vOF5y1YP0eLrxeGwfhFpO8yfB3cJ1dabUW8d++7733XufFixewUkivG/Nriz/eN8vfUfXNanmdCqQC/8kq8PX/q/9PdiE58VQgFUgFUoFUIBVIBVKBVCAV+A9WADoTMIUDGTvwltaA76uAlW2hBwBiZLih+IICJKsAxW/fC2T8CHeaj/e+sxjVaN0JIYOePgnm4UTKU8Ipf1E+vf+4XL31VvngBz/i+265eff9uL9+604ZbGyVzWvXy/bOtTIkB5V9C9l0C3mCoeBHOOJYXvve4lh+eMq34AlnF/UIuoOI8I61eC82EjgJx8yb1jwLiGUb+hOE1fXpgqphmY7l2rz3ewlEi744TLELxNP91NLptZwyFmGSjOrHOra12Gczz2Z+zt+8Ws6nAXbWa+rbNtoDrfz2nWGIjc5NXfuzNN+NRt63wqlW2369fjTiT30u9FyBshUw83n0wbfXfpyn41+7fqXcuHWzhloK0GizmLLu0LHqa0J/KZUuwHXCMruGa+KimwJQ53y/qY9zsV+hmcWQTU/HbBKIXWjBO3RjKjE3J0wUKcStlG0+t7h+i++bfG9SjyhTDoMYDqM+z7OkAqlAKnChQAKyCynyIhVIBVKBVCAVSAVSgVQgFfjmKyBIeLOsEIjARfzS2GQkCPvAkH3qDnhTczoFYMGjBFQyubv/MWF/tjQvmd9TjDmTGWCIdwF8gEcgJEDKtEIq6pug/fnBcXl6cFK2926Vdz/4sKxv7pbr1/fL9pUr5ObaKC9Jfv/owUNOdTwpW1tbZW9vj+drAYRGnPZIh4wNoKM/QYsnNponzCLECSDGOM5hgmttTp6wAGG8Az9Rp8KdAFG4xvTPCbEENrrGoh/6dn1dTons4WSSuwjMPDFT0BRhjlQU4tjekxrtw5Mbve4bAgko6jA3P2rUFDX0nWGUztVQz2be5lgzRtMxkLR+dGABjNS4gqPGKaYGusRqz2rinK3jtx+Lq36zBOhik/zWJWaxrvd+dKz5obuLfuKwAE+TDP5U2xryKCjc3Nks77x3r+zfvEZP9oGmLD9CH3kyO2f/Db1En7V+Jw5ZWGNNPhNOOpYHOsTYq7m4hnDeoZ2nlZq7ztxy7l+jAytluAr8fBYAlM3lGs9g2eL7OusizHK5x/U6nyU503RFvt4MKloareqdr9/81Kf5NxVIBb65CtT/D/LNXV+uLBVIBVKBVCAVSAVSgVQgFUgF3lCggSBvPIpLwYQlXFSQIOoNeLbGI44ZNB1Xl7xOurVkOotwkdkXwOHCuQXqCIeYJ1kKTWYTYBH2sfOJbi464dkCmPGK0x+fvXoFaRuUG3feKsPNnbK1uV12tq+UNjm67n/5sPz03/6bcvDyBYAGSIETaxPHmG6kUxL9E9yIEwkgRafCsYEhfITuhassoBlNVqCnWZffzjfWx1wsXguoDFGkBbmzKiATAE097RFq45yXHMc4GNT2nsRpuwW5tGaArOpwquBKq5xjeBCACfktHUCZGsU133HCJzcCMQFMjAxMUv4FCeeFiZboZzUv+w3gZT/2DbBrtA/QRr3V7vHc/8Src2z68dvwSMdz7k1pGJF9rTq40K3Ovuro+6ZdXNv/qoH3PQ5M8ETSm3dulnfeead8/vmXnGpaZzTgVFFBYBunm2s3stG+PDBgqEOMgYSUM3KudVlb5CwDnMWcmKgATkgmFDV8c2PrnL44zED6Rmn21e8GgKoJmnN45oLt6/Z5vkPafnORPePZU4Dr+eHhq2jPH4by51zBYPMwv1OBVODyKZCA7PLtea44FUgFUoFUIBVIBVKBVOASK3ABOlYaVIyBW6hLaCVkYW6iecDPkDROVJkBDnoAhKFAx+hKEIfmK/7xSsBTYYanC5oTS9JyRuL1cE2RnP7seBynGk5Jnn9yPAKOnZRHzw4ib1hvfaOskfT+zp275d69e2Vz90o5xekFkipdIEoXcDTntMPllDT9uI42yO/VE14BS7q4iIbAK11IG0NOriT3lBBJoCVc8XquMwroEs4nAM1CVxMzjtBJcomF20oXl/W0Sjn7lbPMlaiDfXmS5oCTKAVmi/kggGCnQ54xTEpCGYuuJnNnXYy/gjzVOQZcE6zxj7m77HOmS41nFmUT1Dkmr+K9p0MGFGP+rsF8aOrLJkUb+4jKcVf/CHlYAI9fu8t8E3V5FWuhXRw4gMb0ECXA1WpetORNhWj2J9yr36/dZe67z7EVMp7zJz8brrmtrc1y69YN8pFtc1jCSw4aMD+YudrY094AWMqukbS/BfDqARB76GrfC55N2mPAV9XTnGXhXGN2npApICO6MsJrzUXmfZdDASo0FGx5EIMOQn7DAFgVYFaCSn+/Iz7GBpOPbPmKPHpn5Es7u3//C9eOJHVdIUT+SQVSgUutgP8OzpIKpAKpQCqQCqQCqUAqkAqkApdbAfjMzBMr4QhtQyqHQA3BGMnMl30+DSgBh1TQ4jOLwE1Q4bcfYYh5wsjzFPdCmAbMTEfjcAH1hCmbHDkJdJtPzoFcnbJ37Vq5AmBh8PLd998t7929g3UNSEbesiEAa438XluDTrmyMSh725tlDwjz1o0b5caV3bLL/dbmOidGClMqWNK51czLuTo3v52fkMzrBo4Ir5r1sPZYa3V4VfgjkBGSdYBvJoo31LPPt06mLmOamN9E9VEP4GIfwdsAN47buM7CxQV0mxNKGK4q1meuMnOYRfJ85tFo1eRYizEYV2jkegIKyX/e0DXmzHYEGFs9971rinWt1ifMcz5vlmZ/mBDt3dP63nnYb6OL3w0MtL3vhYHOp6m3hga3bt4oN/dvxDjN74FfT4A77/0PUKyI3OsupD1gVa3tz/4dx3pNvz4XkjnGgvdTflv+vtzHZm5vrokTNHlcf5sMxTkPszP64uSE1ls8f5cxtvxtul9OhWdVTO+ypAKpwKVWIB1kl3r7c/GpQCqQCqQCqUAqkAqkApdVgQuEsBIAAOEjiMjcBP3bZdm5QkLzrWVr3jVxfLwSPAAsBBAdHFhCDHNCCSh4zHPwCt+GWAo0KkQROFUnkGGQ21tEbQKxSmdYXhEytxwfl7/5iz8FlpTy7nsflG1CLDs7G+W//Cf/qOxt9srLZ4/JjDYlnJKQvD4uISCOifCHuI0GuMKu7GyX9WGX8MxtQAoAi+dd+nc1JuC3OL85kAjGxgIFOv5nkPBHN5duK+oBrjAfsb5av0cYY0AY810JpjgGM/KPsRifm1OtgTQ1bJL10ke4vYwbxMekG2se+dhwrakZ/agJTxkdHSPM0jErjFIzYllDuwidZD7NSZXWd97MkgY2YQw/Fiau48wi3mK0uNZ8FmGUrN9WAiZLBYLVAeh95AuzQuyz7e06HkRPzmuJs9ATQHXVWVxLgCnuF65J2MWzvb1rZfeK+fE5lAEHmT+K+aKNW6z+p6f9dgGKID/0EZgxD340M+ZGTGRoKnjzN2b/9il4HHC6qSGWI9yJp7jIrCPo8ndoHjLhmvPk99vqrICg92hmuPA2fa0zqQM+hg2XnZ2d8vTpUy+zpAKpQCoQCiQgyx9CKpAKpAKpQCqQCqQCqUAqkAp4cqWn/0mNtNasAybWgBTE9QlLPKEywAiGpwUZ0AEiVBVg2KRxFgW0Adac4RTTlyPYmJ6fRXvDD/f3r5cl8Or4fFwOT0Zlc7MPHmmVw8dfln/zLw/LJz//y7J/+07ZIvRyC4jyux9+UM6O9gjB45RDQi11ms0mZ9yTr4pJ9qBqQ+qtbwz5HkSIo24j3WPCMecjpHKO1bFVgZKwSf7jc9dgPYEM/5OOsbaVwwzK1gGgNeu0Qg8o0wIKtpDD9bl2E9HbvwBNx5cnMuoWmwOPDMu0W/t1UEFZOKYAP0KkmIt6CpmcbzxnbjjGYjuYYw1dreGIHZ7bn3XbzptPlBif9tw3Jz36XFBoHSFe3SsPIGBe1HdvmVgFe/ZjXR9Fqe4zx3GNxCiu9tl5rsb3GXVdg/2rjRqZK842ajonr9t8PioDaF0fl19f5xZ7Y3gm21SGhuGe15M+hY6Cr6bU+c5CE3VxLgJZIdkQF5kusDf3kDH5Fb+Gatxv8OCOIaW0fzIn5pP6Q59fu3bt/Pnz5+6tv/2YazNufqcCqcDlVOD1v30u5/pz1alAKpAKpAKpQCqQCqQCqUAqANYAIJA/v4VRq2M6esDYYkbOsfFi3pbzyD38ANEqMBIqCDMmkyngAtIRtEXwsSiHh4cRBufTBiIZlmgbE7qfT8aRg2wKpHnFaZYT8kedj6Zl/Oph+ejRZ2UwXC+3btwsm+vD0icEcbjeLetrwDXA08GLaT0ZEaikW2yDfoVYJq43Yb5grK0VbMWN3FwhUZwo6fUK9HR1YwFxTAIvrLEPG2ku080UFMhOeCfk0hqnk0ygZEilY5jLTHBjnwIiQZpQyATywcNsp0OKZ/YdjjFeCLGIZ412kaOMOt3IMVYn3fSJLSs0i/4ljlrC7In2luiXSx1jAS25FscJBcVWvvdd5Iqj6TzCS5nnCl51eB+hnYZ5xhRfg7qL/nmum63F+tV2wf46oiQN4BRz0RUW+dEcC8fcDIiFqMwAvajq/D3V04MLhoTJergBr2NuPuu7J+ztcq5DjT54P5tVWOi9H39H/t5GgDGB5NnJaQCyQX8t+nfP0KVlv6yfWTpwa5uZv8tExszv48Vy+oopblLt9tpg+Hjv2vXjp89wkcXibfAGH1SALKlAKnCpFEhAdqm2OxebCqQCqUAqkAqkAqlAKpAKVAWELAAUiIhQoLME+uikkd2sAzSACMQUBt6QH1Q3kS2FSnKEGtInU6hFCGJSdjHDKQ4xnUMkTS9TAIjv1tfX47sNKNlYH+ACqi4z844ZInh6PiIRO+GaQBjRSq8HGOsYUAgwAcScH59XMAaMsa8+Tq3hkJxjQCPBiZ+at6uO1waWOa5wR4eTkKUDNgkgJEJhgV1Alt/8iW/OINAIFtfx3KWZwJ9n9mWoaWUp4UgKp5SuMPXR8aU2CwiN8xUasXSe0Zg1MA2e881Y9MQz52URjtV5XIzp49UzGnBDTdbp+6jjN/fOSXfYxXPbfa3UvXPPBF3kYCMhvm4wQZbaCtAcI1geU0Whuh7qWGxvabsv7JOPA2LxXKg4p0/XPcDBJ5YyDPLTTz+lIesSfrFHV7a3kHFJOOxmhIjGnMgtZxEm6jAjvpLTQgFnuMgmkw6uwHpSZ7M291d3oIDM0FYhmW6y4SpZv9Av9jggJqOz38DP9mI232JFfX6dE/Sy7DGsUzi6cePG8cHhS/qZYcarJ1nGpPJPKpAKXEoFEpBdym3PRacCqUAqkAqkAqlAKpAKXHYFAnwYowf62NzeXuhaIr9UG3iyAcm5sph3dtFoHZSAySmqwVHa5FcXtjShgKvnwhscP8IM80kJLwyD6w2EO4AZ+na8/hCIQh3ft3jntc/s8/qOQ7XKeEKSfyBO2zxV3b6cpSZlp01/5SJq05dzCscYwG3oCZNwnHBeAXj8bsCV4wNFQEx1zoIqwz2FaZZwP4mFwnrESzqyTsSIRo36R5BkH0IlKZFhhB1cXwRYxngCmTZ5uNqAHl10LfWkjs4rHXahofrwjA5qe+qEZjwyBZzzjHuHty31mXV884exna+T87vOP27qg7h0HOfi/LzWHRfgiJ6a0Ms4gADXGIu+WJPzdczauzK4XtCSlI+iq8sxDVf0u8lnFtpygqhoTej5k5/8v+Xhw8fUK2V7u1/evn0jThttsbc0BYBWx905p5pGmCfj6KwjZT/QzpNSgYt8/E10hIBsJYn3AaZkgSPHnHvruzFhtufn58DWrdDNeQjOQjP+cC/xchvPmBw0sL3G3R5Ow63pcjzmwAXSvbXKW2+9BdD7BVNR3ZDY7yypQCpwCRVIQHYJNz2XnAqkAqlAKpAKpAKpQCqQCqiAMIGkWa0+CdDDnXN61sEkZAjaDm6pdZESVpyWICMglwACkCO0aUokgYcrCCjIABWPj45OygiAsU2opO4w3wV84dt+BBmeYBgFQGKIHcQFgLLgJMqa0J1YTsAOji0ISZ9k/IO+OdYbMIQ7DVAk4BCg2L/wym9dSxZIX32+AkpCopgDHETAYkL4WAtz1lUWvi7cSyIi3VnVOVYhXuiEBra3H/5QvwFWtY5jxxiAIfOQSZpgZfQjcqphjeH6Ynz7sfjaZPVIRL2VpisNfW+Juqv6sQc0dSyL86o91Xpxv6rr/NXTUXSHkf4e6KURjbaSqlXbCL/kOtYVvdZ+rWudgHx8hwY8atZZ86K9XotNzen10UcfxcK2+PW8c+dGuXdnHzfhBHfgnMMbyB82wek11d3Fyv09rX5bYwCoLjV2KcZyj3iEfIbyohG62sZk/xNeNC4yT7Q0fNfC3DyJlanyk2Xt3M+4HMXOt8oV7qezyfQIwZ8tlvMe6cc4NGIXR+Ja6+T0vJEy+so/qUAqcPkUSEB2+fY8V5wKpAKpQCqQCqQCqUAqkAo0CkiTwB8r9xVxk0CEdUIB1wATXMKSoAgLYEvN0QWEMFfWCpgIb4Q2wgifWWwUOaLORqV7daeMzyp3kNV4AqL1Taw/xSlm6eM+mgFQOh1OI3Qc4JKhkIZozlZurh71PUfSvjFkxXidYDzkNPP4S4pupwgTbMDYCrRIaxp41szbb/uKBrqoGCccUsAY6wpOLD5rHFmOYBOdUAHvcDU1a7au64t+WV/AJfqZCauYnnN3fZGc3355bt2AX+ipJsIhoVtFfX7bhpxc1I+6MYg3XtRnb34LxGLWK5AXa2aci72hI0M8WSlduF9802BpfXxw6hHzQQOnPWOdoRGD+Bw+RaHXEAEhmr6pD/7jMIZxefn0WRmdHJf9q5tlc2Ot/IPvvAvQqr+Ply8Oy2w8K6MloZXqje4CTp18mvk8eGGOBpwAwfzq2jGBEYLJvZCVp73eIGCYgMzfkiGWusjMTyb4Q8eW4MyiA475ul09VrLJD3mHkNpTtDxlPd3ZdLpF/Q2g2+jG/q3l6We/4HEoGO3zTyqQClw+BRKQXb49zxWnAqlAKpAKpAKpQCqQCqQCoYDAhNRMAVF07ACfNGStAUa2MTRt4i4aABQsUUfYIszRVdSAF981H2LWJGqR5P6U0ytnQC4hi+F4un+8p3HUtx9YyEVb4UQAkxUAEgR1AWOLVR2BUfQVgCp8XgFuGD7gSXAbwVYzH1YoADIJvmPZ1vsoXAQgsjFwRy4STrigQIZJMijF/F6Wel8dYp02cyIXWaVxdf7OXQ1sJW4yrs82/f6QRP660gBQMXbjmjM8szrcqnarMEraG+ro3GA7Dh39Gnpqn2rSFMd0jOjWeg7LMz+WN/cn8FaAMN1kgiNKuMiatdWubSmIEqM5r6bYpbDOvhtHGc7CeB331He8g5evyAnX5ZCFVvng/ffKjf29sru9WUacUjklv5ynm7ZHJLnjcIWRYZMAMh1/DX6zD+HqoE+uNF2G5BwTiqndiPYoE3spDNMdNwWqTWfjGNvfFxcxb/sRpBKKK+blaM2yw7qu8P0YzU5Y2wKodoN6Uz4PdnZ2jh0L4BZhmdSrIsYK808qkApcFgUSkF2Wnc51pgKpQCqQCqQCqUAqkAqkAijwGntUOSABy7PjozLd2RKAeHolxwK2drvdwTXut2eLaVdYMgNocM9la9kNQCEUqR97lacIUCxj8kuZqL+Fa6rtsZDxfBqQbGJyfuobhqjLx76FKubMahLOd7kXlpmin8GjfkAi+q6wim+IkN0KdJpnEBT+V+FZHTOmE/NynABKNPJaiNLrcC1w8xlExfFaLZLYr/JkeUojjVbthUTVDRWnZEJtFryPtvTn/O3X0iEksAVsowaOuD7Q0JM+gWJOUBfXCqBZtwlVbL7VoHI+5mOfIMtYH/OI+hGKWfX2vS4r5+BHkMRXzGNOdeFVG2fZgjF1wnUY13+YWF1XoDD7AP65vyjgoQJ1vNpvUExXshojVuggUdg/v+l/Afx89uRJWRt2yzvvvF9+9KPfLfv7+2Vt0Of503L//gMmBBRDmxGhs6I9whzDQSac7ZPk/xQo1m31whkmkBP6eXKmytluyhjuQSdOIAWMMWeB2nxBeCYcjKNY43eDI3HZafUjzLLX7cPJlpuMtsuedxnrmNDaGcB1n5mTU2/6ij6Pb926U7744gsO9pTiMmSWVCAVuHQKJCC7dFueC04FUoFUIBVIBVKBVCAVSAUuFKi+pAZ+tFobrXZ3B/i0I1SgVpxkKcCoEAy8sljCklZwCrDSA7zoRNPRE2CFrFokgirHJ2cBvEzyLnwyDE5XkIDDEoCK8MpIGC+8WQEg6YRgRAMVSItwxgpqdDU1c3AcfU4W674Jv8QpwiLBjfUM5fO++XZc814FhaKO/UYyezoSHukkCzed62Fe1mcAh4oSa0QOw0Gj/9V44RBjnLoMZr4KLRSStVrICBxyHvYl1LKoRUCweEYV10wHMa59+ZxPaEh95+oxoxWmVbhoP67fNTmfWB/3sD/0B1zxXLfaUmJHsT1Z5ZgL70Nsvv0VUKIfbX2Upp8G+lmjufad6yQ9XWjFReztO+99q9x763a5fedm2dzaKRuba2V8ehbQyrauVwCpxg45HA5LdzEJXQyXNLzScNs6j/Xo0xxjAtTp1AEBaVzaoUwZAAAgAElEQVTr9hpPOPmSIsS0zoA8ZO5fU+yj7ntkeBsw9g7z3kGjDYKGT4GGA+qeA3AH9rG9vR2/0TFhoFlSgVTgciqQgOxy7nuuOhVIBVKBVCAVuPgPnfgPttQjFUgFLo0CcJGvl6VJ+smR1QdebPBy2DLOT35CCYJm0vrKV4AriyWnS7amuHcswh7DGPUERVJ9yIv/Xnn0+BmhllzzXMgTObhoMzDnGI4qTyi0VGgk/Kkwy2eCnoAkgJfWEtcW7QVAmqcqv6lwqIEu9iEoi8J1tGdkS4UtorYKfcKRBhiyjSAs5mVFMurHXLgMXsR7QZCJ9YVK5gjzfUAs58OHtzyrc2m+fd704zzomJkI2bjGOSVZat7HsFHHMYV+ztf1Uo1xBWGLeM4DvtXR/qOYl0v2w5xijdZ1vqv3hoGGJuhmvi7HpAbb6KxrvTYuvTi9k3e+VyWqr/pbrSPeOS7PeRkHGvhsBS4NbVxC44bLtfKd3/kwxvDESZPpz8ajcIOdnXmQpDCLvGHTeVnb2Cx337tTdm/fLf/r//5/lNPxtJwpOr8N3YNz5l73xp8hvy3mb1FPD3Qwhx1xkuEe6wFdDbVc8C2EHQwGrgU0yJzpEx0UjDz/HU952AfE3sE/NsERd8yejdGrRyhsr0ssbJgWHShLKpAKXEoF/Dd2llQgFUgFUoFUIBW4ZAo0/wF1yZady00FUoFfVkCKRM55qANuMbiCZcztWMjgM6CLIWoBLPzmnXWiJ7+FNrW5KINTJAEjU0DKEc4hg9V8J+jRZea1fVhsG+0Jl2uuhUNNX+GUos5qzFqXESzWefNTnUmv59GMEZX5Y/8+M8yRlnHvO5/5acIHBUy6tOKba4tt3yzmwYpnACK/HbuZs9+uUzBlH01pxvSAA+u/2aap43fTz9ffOyeL41X3WNz+0p9mrrFWmsT3G21t4FoFcM3amzbRt/3zad41A8Q7ydmqOD/r+G14peCsw74P1oalx6dNWOkUYDUm/5quQeEfFDWS8O9evVK+9Z0Pyu//4T8qLw5elc8fPCxTujbA0wx44ShkHEMnxybuZ5wW7bvCM6Eb/TluM2/rT3CTTSaE7lJXmOY79Rey+aF0eWduvV2ur3Kte4wzMtuco7Bcp66OyT79ushmoV/deF5kSQVSgW+2Aukg+2bvb64uFUgFUoFUIBVIBVKBVCAV+KoCzX/2NxgAZHJ6ety6srhmvTGw4Gi6XI4AX0OAwhbPBGRYyQKOteEhEASSzodDh2thiy1hIC0dSdQzBO7VAXnNqMwRglFgR0ALqnGBaScAhtzEfgzVE2jYLgAHHRr+p7sr3tOPYIqpAkkAUoYvAl86HilAccyvF5/5MZfZhbuMSg1YsW9uoo5zuuA/zCXAjx4k3jt+nPRIaCA0sAIq+hV6LXCdCYiEMLqmvjIPx2dNOuxcm32F68p18D8BoMUTQi2+j/GEP/GPIEtRdegJBK1f11Q1rJDIMWvbqoF7s9qRWHejjMn5zfkV86BGuNFwoDFKPIvTEKzs9JyrvdA3f7jyAIeqtSdKup4IKQVGmYfN8rpNxXmcEhnuMc2I65tbpTPcKJu7u+X2OyTvv/1Wefjl/fInP/mTcjYmj5jDsFYBJnn1A4LNujW/mH1HeO6SXGNz5sX8XP+AAxCWF2GW8wizNGTTebhPTNKmSxhb6a3HWRPA3tmANQnC2qxhye+tC1zb4BkHUrTOAbTUjkIHWVKBVOCyKcC/cbOkAqlAKpAKpAKpwGVTwP/oaT6Xbe253lQgFXitQMAEbue4cuYTEp3DfXimu2aD7w0ggvcBJN507fjvD4vfDfwJqMSzps+Tk9MyAZ6YqL+pa52mnm4g8ZMww2shiH01/27SUWT+LOFTBULmMeNEQwEbwwu4GsdZM+ZFW9p4HRDHea6givWduQ6qlbMo5uafZh329WZ/FxWiEv/uBIhFXToibC9ee3rnm1r4sM6l1vXa0vTdrCce8ucr96zZ+rHGFSiz3pt9NO2aZxH2KNRajSPtexMKxsmVPBOKRUGAi7pNZ3w7v+Z5o0fzunlunTfna70FIbN+W6xnPrFZADlylAm+cH9dv3WDEMzvlzt338YZNi9/8rM/L7948Kgcny8KjOxiXPteMj/3R1jqoQHzWXWrNfviOMJU763nRw0iYT/X9mFhLkTItlv+vnGeAXpba91O7wrvr9B2nXaEFcfvXYIGs0wuFsLln1TgkiqQDrJLuvG57FQgFUgFUoFUIBVIBVKBS6qAeauiVBjFJQcwBlAx69UWiITT/bSTtbsVfgAaSAImO7FZ1OWmmpuAJZFAnWg1+EiXcEkdSWTtKgdHR+HqaeEcgmRUaAFc8pTGBrAEDIlITvrFpWT4IEFvXAuJBEfVPSXQMmwPTBKhdk6mgRmeZNhtA9cKSd6Zn/4p+/UjvtJBFoV126YZ22fCLkP/LCayr/3SyrG5d60RMkk73WC+Nz8WF9xXLZxohC0CYcKGtoIzb47jI8MEG4gUA4ZVS61oFmGDqzUxtim3Ot1B7Y735jcTGrVwztU5WleN+KCRWkGJ4p2XTC/mJCAkwNGRolRgSF8+s5LFdaia/cWD6niL9fMuRIzn/l6cS/3Y3mvXaTSuOnlvvjOBlXBzynXs4bBfhiTRt97Z6SlhlU/Kzz/6vDw8nJRItc9UBKcCR38fJCKLtibfH41GAcP67JPOQXYp9ni4NigjHGTTOTAO/axn/rFeb+jiY8YBM5dz0FdXsRCobM2W83vo9pLxHrMfbF1EGENeW/x8K/CMxrEzXilCllQgFbgMCjT/3/EyrDXXmAqkAqlAKpAKpAKpQCqQCqQCVQHpiB+zjvnpAAq2+VzjegPo4Tux2Jt0IEBabS4kqRDCe8GPLjC/fS4I0UUkPCNB1QWUqjCluoFsR/8BeARgcU3b6jLTXQasMKwPMBKhluTvcox436vf9hdOtAb2rPq07zo/gBjtmEAFSa5qVRzP8uZ3Mwfbupbm07iUBDGxRtcJOBESeq/7bsZnwQmMSw8vIC+Webn8jo8Deb2CLbIaoVSjoeuwOI7F8MsKmQRoOOwaeEeXzRJsay+CsjeLz6PfAF60X71ucXEx3oVedvjmFtMT8240MbQz1rEaIPpmDa49tMHdZV3n32FPLDoBvfe5wMoQy4nwkH00J9mz5y/Lv/7Tn5a/vY97jOGJmvwKNG3GdqwmD5m6T1fa9AYerFr3TRcZUkZxPtZ3/v5G/AUzz0jZRmilKvBZrNP/LQ4nuMG97jHnu8b1Nm2H/paypAKpwOVVIP8NcHn3PleeCqQCqUAqkAqkAqlAKnApFQgg8pqzwA0ACrpnIuwMSUadVvcQKDGFqAS5AVZYBB8YoVasgVc6p6BmAanG8zGHEOL8AVIIHgQ8ASwKIZZQDKGFCdUbAKL0PqNi7QcYNiMkU0eUFKhDXwGOdA4JYHCJ2bZtXjLutVmBfEobXhIACzbiHP3U+EKcUPRjqF8XSGabaM93eMuYv6c4hmtJyiLMoyiMzMnQvpYgbNVfnPYYFXhOH87TcZUjEsRPhTiEqepy65GQvsO5nkwzxqX/4Fi0EXn5LPpdjeW8dKjpYnNdbXWxYydDsW57Fc4pCHL8cNX53QCt1dqta7Pof0WPHDX6YXw1a1X7G/VW6+OlJ2LO6DuKfaKNbrAW4zp3+xOYcVGrANacLkdY1nfOuSM4A4axnj5wbDI+L+c4xg4PX5Wjk7Py6ui8/PTnvyj/95/+VXlGtSkTdbau3/BZXXYt5whgneNIm6PBCBfZOadhtts1v5i6h5OOuQq0/ASkFKIBZec9f2Oshz/qbN41f2ABzToBgvv0zYEUJupfrLfbPYbnHNZWa5N6pszjl+QqVfh1aW7q6l8/z6tUIBX45iiQgOybs5e5klQgFUgFUoFUIBVIBVKBVODvq8BX/jsfyDAEIEAJ2guAESf7zWEOpI8HQshDArqsgIMDREjeaqTmnZBDYGSK+dlsDLTgNEtgWQUTnTIHIFnHe9vUvivQ8rnPdARFH6u8ZbqOfKcLTGdSjCWkoTSQKYAMMKXpt87n9ZyDMgldJBz8iXEBL2CR6MN2Qqum2N5/agFkLcyvVUMGnQv/C9wkZiM5FsYwQB1gbHR+VhZkhNes1B90+azVteOsas+FcQAk+ZOJ/YFxJv5vG5LKdwMOa/8VxTiPmjPMRswR0NOORPnuCXWYSNWKflfFfQkthWhB5FhyONeaGhWI1RFW1/QTa2Y8nWuOFlrxbV+W5tt6QjI1ZGcCPqJIHZN3XHLdCeeY7ZbLYYQ/Giq5tbVVjkeL8rO/+dvyEjim8QuLIk3IS9fAv9DdMFL3t+6VaxSS9cljNhj0QlP3bDoRQBqS6UgVOjqvOful427FdmNtVkBln3Eo5nLCekgb19qbTObHvDrl3kjP4cpNFlPjvvkRcJklFUgFLoMCCcguwy7nGlOBVCAVSAVSgVQgFUgFUoGvKtD8xz+Epj0EXhheBu3RWlS2ADfXSAY21J0kvBAG2UBAErAEt1Fz7b1gQk7htVGZA2BGD4jR1f1FQ+tamu+oR74nn4aDi1Frf8CRri6i6hLTHRTjAUsEYgGzIlqOhoAfYc2UIxDtR5BiH84Fo1A4zVaTwpRFHfkU//WjA6nTZbYdWnE9Z8kRh7ean7m+nG7M1fUKsEgqbx4wIVeFQ8wLh1WFdBWSBSzDwTQZTcr0HOfa2qR4qmJ7BiBTC0IDI4cWcxOkCb9iHKYSrinHN9xRPf9/9t6z3bLjOtCrk8+5sXNAzkyCKFIkQYFiksQRpZE1Hj8zemyPx8/MF3/1L7A/+7c4je2Z0SjLQSIpMUikSIIE0Aidu2/fnE4+ft9VZ99uQAAIiQDZ3ajq3neniqv23t3rvWutYkS2OwvIFTZWIQchTxAhhW1Wxq+7psn+KSv7HVtArDwn5tFCzOsWVWJ5z32ucwPZgteQYdxgvh0nDXCqdKt66IF10I4utDE39Fk5WOs04pCZn3LMvc/B6nEeJe53eovpxs4gvXZ9l2hx5uZZoW1XJdUVk+FGOZ818GzMoX0YAVsnk27Es2vybIQ5GzkN4B9zjWztN6exDfsjnj1kzfxElcglxo14OB/S/UOgmgHRHud50o34ZTZM/3AGbTV75BGWvXk1S4qVVCRQJHC/S6AAsvt9hsv4igSKBIoEigSKBN4DCYQSRD0qGSUVCRQJ3D8S8N1uNFvNxcXFDkhjCUhgDLJzgIcTvO9tYdEY+MA14ILvf4ZCSsC4UH4T3AQV5hNg6RrnuW6HU6zGhFwDLIdM3rec7Wrlo/ujwAfbNe7mLeJecb8CYpCOyC+DsV5jWklCws0QSCbCsU3zB+CZ12Ne67Sc7QnGwmKLdr0efReGkUHLLM/JxiizFRY3uMbqnlSTARDQaG6VZX0SHU/bbQDYYi/tMl6CwaeD0R5jJHB8/zD12620uLyUWm3cA0VCs1bE41IOjgOpMSbH7xiVbwZT1u+46AAWYIyZfKAkuiQEY8+fyuXSUo5V669qPrgUYJI783pjYF6mTmVODYohplSA5JwhJ4PUe8B1XSurZL1VqtrQHTRkPgdQWX5AL+bS/tjrNuNaXFqJOd/d30sbW9tpTFdEegHI6HPEEVP2eaKimZD3vEnrCkg2ty7UktCtmm9lZ547++i5br32RVlyXvO5qzebU/JPAY9dnrtzs9nogAZvsDUp3wZouoKrkokUz80dY6+ul32RQJHA/SmBAsjuz3ktoyoSKBIoEigSKBJ4TyVwp+LxnlZcKisSKBL4OUgg9P9MeOBcAIrDbnfhNFZGD4ATHsUN7RhgAPzRgCkJUrIrn7xGYABNij4ffRc8D8gFCCNW1Ai3w4ZwApOtKh6ZYCriWVFe2GNZ64rg88Qak0mAieKa4MN7wiaPdT8MgAZICnACerFPWoVFPi3RtDLC5S6vpJjJSs4L76F7lg8LKk/CYgrchJWRwf8FM1QVPRCsCHYES7ruuVXAJ/oVICfHRtMFUPhHD7FkI99kJW0TqL/F9REWYnuHrKrYpX5WWWzDXaaTJdxMWSyx3SE+mXAJqzLKC3h0s2Qwsc2Af44ggJkQqsYKnbQ7wY2TSFq0R2O0MdPay0T/nVFjwZGBLf7GLc+r6wI6k7VrsUa3o8nIQ9uOdUqdoLfIx+lRinnnLM8bB9y0trDa49j7sSAD1+q4lArGnPPRaICl1ywdDIZA0lHa2d5LAy29yOeKpzVXJmVObLsJpKRj0Qa3qZ8xC0Dj2TEA/yANeVZcDIARkA93Sp812hJ+YXIXm8+c0K1a8VKjSPvH6pVI0odL2zJoo76gqd6l7Cp1rOIau7m0wPoU1h1/8njtS0lFAkUCHwwJFED2wZjnMsoigSKBIoEigSKB90QCdypJ70mFpZIigSKBn5cEYASyk9kUSGNQcqL0N45xvoxbped7bFCHDAkACDPBF/f5DFiU6+wEJkIlQUkGUhkaTQFF/T6wbB6w33vhPii8EdpQh1u+noGTgMxzgUe0AUCy7oBYWldZJtrlpzDE2F/UpbVWlSzHAgNkrcpmUCNkgZhE/d7z3DheYLBcp+OgLKML4BQEx1hhBqAXZgFmhG9Cq+gzDTaxDmtx3VqIZ5VmjLW30En7OxQDZo2G/XClnADLugsulEiXBWiL1IHrYY1w8BMs1PIYgWWM1/hZwq8sF4ZpGQCPJlcRw8yOMXbhYwV+XEjAcQvRrCvilnGshZsVKCPTkdyjVm45Vo61khNZKRevzbNb5ChVdXjhzmPnShnaX/sXdXIMVYy5Pzg4IMA+cdmY2y2C9F9bWyOPrYIVbZ7nRgBpPdbhDE+Ff3TCzevCQwEY9oxHz5rtaEXmdct7HLHgqFTX13BPnQ8kj/NoKC3K9KjXuGOHlOvz7LZ5Tldov8d5fXX1eNra3jgq4IF13DnuN9wsJ0UCRQL3jQQKILtvprIMpEigSKBIoEigSOD9k8CdCkZREt4/OZeaiwR+NhIAssA5qrYWFhaagJ+WQc1hCn1YwA6gZR/gAisDVAhZ+Mt3QKQRsEAQEysO5iteZROUAH2oXgA1waprY30zIMfQGFhwE10urSaqqmCTcEU4AtjQ1bGBVRXVU057H2JLAcLsRAVNhFRaD5kmwDFdEN1M9iv2Y5AMlkZV0kqpSeD8AFNH7Qu3NCIySHy2mgqLKC3W6AMGR/QzGCF7JGDMMsoagD+ADpULxoRLdWJjjQkkbzyzOKc++w06xGBJe6TsdtpbXmGclG/lcYWVE23VhD3NDA4bUy3aJliX5VhcdQCQc2AK8KOA57LTKs8+uSkfs8kOncgAaUIyj+OSfcjgKS5grWV55ywC2guXwoov5488d/yYTz9NzdtijNGmc8646Sbz5zziRkp8slu3bsG/Rml7dye9+vqltLGxk9a3DwgChoQEX7RG0bAGDItA5s7nwPhxk3ChzauaMrnIchwwzPl1jgRiTazEGoKzGJ9z5XionCkVKta5ftQ/liS1bso22XfYT1vN9tZkPNlmPDUg8SLXWA91Vj95+lR9a2fzSG6KILdxhzDKYZFAkcB9KYHb/2rcl8MrgyoSKBIoEigSKBIoEngvJBBKxlwpei/qK3UUCRQJ3BUSkITAZlodOAUB+acdWEGLPaAgtbFECmokEDHpDpgB1BxwxVVhWAZcEyyoPB4BMQQaNSzOtre3w91N6kbhgCvmMQVMietaVAFGAFXGvbKNsPgij8e27zcogv0DmnRB1G0wVq8kj8DEbawLIn/AXXbqqC1XwBRoVS6bwpUaAM/hGX+MA2rNiRhVNKolE32gy8b7gpTFTWGYfRG8UZJA8DkfudJkQNvmJ/i/cMZ+61ZpnC4Bmal/cEj8sWlaprFmt5e6SN2g9lGLfaCMUGtGH5TR1H4gD8ceE0X9Bq8HxdFFxiPs4lqunhzko/OUUb7IK0aR+277UQ95qvn0/M0p5BzymMMljr1WzYFgspo/yyoLLci0Ynvpwmtp7dZGWj52PB3DCuuwf5CuX7+eXnvttbS1u59ev3wzvfDalYQPKrJljuwh7rEBG+nzTBBKoknaUB6cs4UFGVZu9kPwpvuksvJ5dC61VIznbpTlbn0hy6gtj5v+w1DjWdJqsk3+Mecb7PdxvV3g+BTHy95bWlrqAY2n+/v7miZWj8a8trIrEigSuJ8lUADZ/Ty7ZWxFAkUCRQJFAkUC76EEVE5KKhIoErjnJQB+CN4SLzRQoN5utYRjS0CLFUDTaZiAQfpPAqmEZAEzgCB1jHAAMhlCcP8N4ESpVODFe9Xx2sY6AAQgBRCZAjkCtJCXZi1C0j1OyEKnsGAKKKVlEV0UhAl5OKJLxKICNo0BTAKUIe6LpjHue+YIN0PapVMAJuHSSCMr8upKmQGPbYbFFv3RYkk4EzBJeEal0Tfyms+A99Zpn1vAKFOAHA7Np+GYfbS9CStc2pbuk6NhXk1R0NbqCKlmsZKlAG9EPvf7WFS1AD2px6IGxCObMbYkk6RdgY+umS1WvFSOjSZWUlTOqMMFVHfCsJZznAqCpOzscz7jRFdQrob1H/kiAbboefTT6yYhY5SZ75FamtCWd2NlS+rPsjM3ebnhHGB1FTKwj2FFSLk94N9/+A9/lP6vP/jL1Fyop/Pnz6fPP/+ZdPbUSVwsp+ni9fX0Ny+9nm7s9hnzAmNT3tm1Mqz16EPV3xhJ9COPw5U8dSc13lit1iGmGXPCHOKUGZCsmjclgXijHselTJShewcFcNMKMsYEXBsyFzvM6Yj7J3CxXOTeKxx3WvXWwunTZ2f7+69I7BRcSUUCRQIfEAkUQPYBmegyzCKBIoEigSKBIoEigSKBIoEigbkE5AdBSQAyxFNvGJT/GNZMXfYEy6qdJHj+SSx32qCjnJGLWC/BS7TsEVLdBkpCFC2LKhDlPSvX1un1S5cD+ghXvE6mbM2l9ROQqloJkUqBVbnOADfkE00I5Kw72qNMDWuuKaDEPmSLo2xVFLGorN8EJWFhTmCO9c3by/5/WJHhvkfvhCbCMSGZoMnjys0yV6LFnKNno10XK4g2jebP+QhIMx5jNcZ+Soyx0eEBscd20h5xtuhZDsoPJGtgUWYdzYYunwban8dNA6Ydzg5S24UGpgA7oFan1zaQPH1rBmwT5lUprKKS0C9b6ym7CZDJ65GEYjFe58fA9hkOhcwVPn+r5DyZlE/MJcf5Gn1lbJF0J0X+zkmMmzItXEM9lheK1qxG90/bqAOsXr96lf6ntH8wTTdevJJevvjv0sljy9GX7f447U0AVe0eJZkb6hdw2X9jl02Qh31WnhMqiWdK91T6np+tWliP9Xq9uOd8LywsRn8ODw+jy1GeTiljQaP7Sj5xT1zJfS3P7DNjmXAdTlfr+B5wb4ltkbk4WF1dHbGiZV3rtDvS0Xtzx7VyWCRQJHAfSaAAsvtoMstQigSKBIoEigSKBN69BCrrjbf+5fhczbxTp3r3Vb+LnCqAKipaV7g/SqEMvUGXO7pVDooEigTeWwkYZP7s2bMs21c/BfSJ4PyAg8MW0GBWn7G637SRYZJgSzCT4YO9EDjwA9gh+MqARXhikHldEeEXWDzV06uvXUxbgKNOp5OGwJcIdK9PIJBFgAGRAVTklQqrLwGraVI+gyLxkqs1ak0mFMlB/8nJ+dAVM1nZ0HZNTaytrEM4EvBN+EIfBSJuwpLbgeiBXACYOsCvqRsl8MdxCE4cUyTqDbZEX4bEOjOe1uHBXtrf3E79/f2oU1g0BZRFLDTy+T1bWFgCcA2wVgPGIKawoAsLKOCegInvn3u7PRwcMhRWXZywuqVEyv52BVXzb7NwTlkjywBFykxwRr91U5yFRV10nC4DzQRl5A+Z0Bf7U31jq70NByCaf3vFgGFVxrltzeER9VMPAnWW9Yi0vPdmnAjXTF6LGGmAtH2s+WYtuRp9Awz2KX9pC2s45mPqmOvGlKM8Q8PHkefDyqmHPtvfNgseMPoAYRHzzbFTlzLxWfHZGrMiaGPEnM2t+qzb4xFVOb/WM6FP+E+Gi6/1BwikUVdMHfHcKLsRschgqD1WyRzyZB8wjjpwsMctYfFuu9nafuqJJ2cvvPDCPK5cDLf8KBIoErjPJVAA2X0+wWV4RQJFAkUCRQJFAnejBEJ5o2OobvHnDpUUBcwea52gqpsVVvfVucclFQkUCfx0EhB0CBcWl5d6tUltFaunBVCCAAOXs8aMlSGl6ARu4mcDjBTMhnUePcgv6Rs6ENcBX9QgqYjlLwVk69u7xKC6lD782INp1B/4QgM7soWTXwCPO82u/IfE9wAQogVZRm/5vRekC9F0YQTlhOWWYMx4VEIzvw25T+OIT2VNQh+vCUd0URSimC+gnFAG4NfwGyOkIdUdqJ1g75WAQuxHtDnuH6aD/d10ABzb3dpOu5ubMKpGtNWBshi0X+jVADiGpRmx2ISPUYd9sNcAmzpjiO8YjMbzamEB2+9jBeVYGtjstQBDwp5eL4SSZkPGjgWavQqLKGKTCbKmyCrgmfKJYeQxH31faaNK1ZzdllXug9cDqrE3hdw59rp5Ay4xrx7bX6+HWyp5jYeWYd00DbCim0KXZmiX06lWehA1oKMzOcK6bIJs7bsB+G3JPuY553g+Dq0Jo02GbZ+qvlZ9UT7On+eW9zyDz7mbLkLQwtE8uZ5cn+c+6+7dGoBL+tJjqldw39xBhut0qYtl4gqPwwMcb1L++tLSSjp27Fha33zjipbcL6lIoEjgPpVAAWT36cSWYRUJFAkUCRQJFAm8swRuK05vlS+rjG91591ey4odqs/bFMiKllYLlfKjtYL6qgk1J/aoVKq51IJGOb+S929X7zxb2RUJFAm8kwTQ/0EXhB9jj7mVryG2VY1Gh9ewh+dem1Nu12rtZhPbGtDOhOhUHFnOIPhRfv6e+poH3PB9lXoAVKgj8oAz0nf+5u/SR598Aksc0cgctmghxr+MY+8AACAASURBVKlujRPjcQFPDJwvRDEou/Xr7geoC6shiF1cG+vOCIASkAlIRqyUaRKA1GZAGToTq0baTz4j1iMUsUynaR5Xj6R+45QZOwwiMrY9oI5JwGXyyzNjxU0twcaAvYh1Rr5et5tWHnk4+iacESBFwjLJr579wr+SdgExjM3xOqawfKO8fRH0qYQJ+JpAJC2otE4T+kwOtTKjH5QVjNUBcK0e1mW0hcsfABGXTmtlXI7ZMmDL2DNn0Ra34/7tvWPiS8ouemsFnBhnLb7RcS4fzECpmtYAe7RjoZAKE5ZrssAc1nFkX3b2dvlKxzNF1YJJIR4rmbKPeQVQKi9O6D9yoIxjsexgHufN/mvlRUG6xb1YIdS2MxDUgs7xVklrRJ816w05IN/p1OfB2cvzaZ1a2hF+LB7y5hyUITt9PY/Tn2sU2OJ8uT+ZHOOZepg+XWUF0YYrcy6vHqsDyGL4VbtlXyRQJHD/SqAAsvt3bsvIigSKBIoEigSKBN4vCahVhZ4131fKg/vqmMPbigwnfy+pGJnch5qGMiIMQ206yuux9++8dnSzHBQJFAn8YyRQvWBN4AE2SrUGoPqQ4z54AVhWWwEaLeBwBkIK66IZLpPghUYNN0lXAoQ+ZOse301BjpBI8GOq3us24GcgiOLad777/fSv/6vfS3VWHxwPsvWY8KtJ/KooJ6gBfOCBR28yhLGeMfBLizLoRgAQj7UkmwCh3MZALyGGgEkI5QqS9jncOOEjAhUtxbjAXyzBwu0RUANw0jQuoMqEtv3GTHHdo+yYY88NCh8gjfaEaF2C6XfaqE6LizFOV1hsCtwYBwVwsSQfh405gBHcWE+ALvbNCCqf42jVK0gDcBLgDA4JXI8sHJvQbMa4HNO4kVdsdIzdhV4aDQYBg8JNVKsuZUN5xxtujvZ7DpCUn3W7VXNS7Z2vO7+pVd5qHwOc/7C8VcqtCEEX43G81WINPBYxzt3d3WjbFUOdQyGZfpkBTOeAyxU5eViQmfOS+2ebQrGYP9qSjfm02S4/Yj/mXDkGEGXe8YKMtnx2vC4o9J5zEuOl7/mei7Ha1O36XGAgQF2qE2tvepJ7S5TdoBxdaJxA/q5meZwFKXrMYfP48ePja9c6swGyJ9GpkooEigTuZwkUQHY/z24ZW5FAkUCRQJFAkcB7KIFQWKhPZWOeKmXBPRoPWpNHKqQ/AY6RYZ7Ma0GLkyhv9bfbml/Pd/n55vOjG+WgSKBI4J0lUL2v1QvcaNZbBOXHAXE22qfoAY6UMKv6wmQ2aQFrsMcScIS157QlfCIIGZZQUAvQAS+qKxHG98BA7UCQbJGF1x3AYxxgJUPvVy5fTlfW1tISrohaD8VLzh5CF4BDMKR7HstkAl78CPCmAzzMZ9D2IXDCOF8BPwBdrmApSDI4u/BKq66wPGIQ1bdDWOWxLpzCJ4haqhGoamqQLMZkYHhdImdYpGlqJgDSqims1gBUWoAZEN8VLLWsqrfZkjHOgHT2S19CGjGIfY77la3quAWwYQVKrKICXEl8SNozKSsD3QvPjDs2HXcjOP1YkAfkGgwAcb3FsJizL1rhHQL1moAfgU8bwNjpdZPOmypxwiHdHHGJDWAkEPQaHWPLSWAWPbBjJHfUzDXmLrIxnYxBu65pfLvNFFmPflhHBl35RpwrU1KW8SQJyI4S9TQYp5ZjMwTrQgh1zgVTthmWYMiXTkcR4Zguq7I2u6QlmmO3s9bvpuzcnHdh1dLSEvMF7ALIWa+QzHmwLoGi82Ty3AGRl0c5W6J5neemS3UnqdvFKS5juzdotpsTrPS6POPLZFnE6gxP2dbsIx/6cPre975HLXMZWkFJRQJFAvelBAoguy+ntQyqSKBIoEigSKBI4L2VgApKlThGT0G1+PsJ/5zQA80c6s0dWczvpkZUHd9xOx9W1Vb7v5ehXCgSKBJ4ryRQA7g0AS+80jV4Fim5guXU+OmHeFPugiUgHXVi9hO/HNwzjxEF9zEkutzCYPzZIqyyXBLkCJUENRXkWNveTldu3Eyf/NgzaWewBxfxQ3HbCs2yvvNjqrV8ZiMZjuh6qAVZgClcIm3Pzes6X/s1sYxAq0mb9ikCztNBr9sP3Rv5gX1cKzWs3/pwXXTvSpGuihlB1ig7EsQJ6+IrRTvmoQ77VwPEWJfQRcikK6jJewGbKC8Ki3EDbhrzVSjtkx3NX00/ga5gIDQCxHGrU2c1Rtq1nO2O+7hnwvFGBr2nkO3rlum+wdibLp0gCHLcjlchkGwn+jnfe03ZRn/tY2xm5DplJJ20aK6AUrqEhvyir9TJbdmd5SP/m+oHFQIdKQso3N7aRXZY0THmGgwVwUad1tfgWCAZcshCyPKlPcegJaHPVhubxTf3f4ZQBGpRdj4eg/Wbj4lGbhMWRVg4mhfh2BTXVOuNupkzy0b++TPLsYnHpS4IW2V8XYDkEMu2GbCtAYDrcb9DuZpArt3uNohF1tjc2mTi5sLmoKQigSKB+08CBZDdf3NaRlQkUCRQJFAkUCTwnkvAwMcmCVgkFI47k9Ya84RuOTP2tRnmpUKjUCt0M93OfXQp3zj6iUUDGs0bch7dKwdFAkUC74EEsI5qwgBAE6CpFkBgiQhjK0AgvA/Hm7ABqdMC+xZwBLpSH82hAeGwYhXaKaQMcEYELF5VAUcEZteiit7VdD/0O4Ed2iEA6i++8Y302U/8QrhjDgEpAT0AJMb8ur2qo26K9gggJNQiVeCNtuNci7JAQoCfDOeyFZoWRAIkk7AsuwNyLHzDRc8k0JkBVKZAD6HPRGgD0GkAyxxTTgAfXENtV2uygEMce99YafZjMree8tgxCo+ibfruvtpcvVJbrRaB9ydalHHfvo2BYQ37SNstVm6sAb+mQ/uBCyoWY23ENvEaglQOQhphT7vbiTFPmRHPa/RD8OToqr44BmWb95UFVZChuOaUCBBbjp868kV/ZghG4dtydGzMMIOk0lyH4w04iUWY82b7u8Qf2waCDgFTWgIK+tgxt8yHdShLWGsuS5tzsGj7MW88A8rX6Ytx0BelGuWwXIw/9oHkNSHlcMTqmP5h3r2mxVq9ybPBs2b8MeWOQVnMjbVlyBflCW0Wz4k/nPQuHe1hPclCqY6df8CAZMicKSJuXadT5znrHj9+srGxtakrcrwOlMsdCslwVlKRQJHAfSGB6l+C+2IwZRBFAkUCRQJFAkUCRQLvvQTmagkqhyqUUWXYzfA1wvDBS9xXy+qzHbIN0a9Cc1BFc5urYKE0qTXxV/es6v8g3jZb1mA5OEqhlP39y0f3y0GRQJHATyUBXfaAFE2YVg/Ff4ltgXfTtA90AJrV8HTE8a422QbGsKxl7SQNYmgDBsHqDOjQBB54HmBDMCT0EMAcWQxRQLObv/jGX6X//r/7txqkAUOAX0Ai89bnVkO6WeqSyGIAGFcBOKjzKMEkhBwjgIVQjP7lsnRcsJLhioAkWwu5YqWuh9YfCRhFf+NwCvezavMIZIRMwhOBTpSjzFH9tOmYzGMbAXZoU6Cm5ZbAy3q9L6ixQoTFVxFw1cQdEyhkbLCwKGMEunrOAIa2VeMTONHlj3JEISN/K1aybMxwo6ROI15NWCTAFP0FFOlauEDb9BCmI4TiByn6EP3J30vPHcNbJeXqfV043y7FfNIAVDTGVtWlLKpjy1bHhweD1O8DHelbo+HCBkCqOojKfzSUlzK0zblsLSdU1d1UWNXiGQBEhVWZiy40kR0xwCiTre4sW0FH++YzYF0dgKLA1HPvR7+p2zkQjFbzr3soVUDA4pmK59X+Uy/h2Gpaii1yNETefeqY4e5Z4xlcmBKLD1DmVNR06Vzo9uqHrGg6T28vwCpH2RcJFAnccxKo/nN6z3W8dLhIoEigSKBIoEigSOD9l4DqlzpOi4PFRrP265/5bOux8+dXHz5/9hza7NnF7uIiFhB9Vvy6PpwMX0fx2bp27Vra3NlM3/7B99M3X7yctANRLcmbjkmhG8Wv8KmWENmGy36jrqHyVClfFC2pSKBI4D2UQMYqYJvatIm7WqchKdNAFOsZYA+2NIRTx/xpNJoQ3qrR53gd/jAaT9MStGOhoZEoZkpAh2A0EaB+DkDspqBCqCE0GmjxBRG6eHUtvfCjF9PTD51PgyGQgfthJTbBiorYZAKOHMvL5QC03Mq9FH5EXDCAiMDDunVDNOaYVmoBTrDUqgCK3w3bNhD9GOAm2BIsxX14mXv7pXWQXzfjm/l1sl7dGC0/xnQroBvoyrzG/SJifhwTtz1cHwU/tqMA2k08U0m6lgpnWq1OQDC5v79RMHldsGW8LyGhX71mDagGvNNaTPjmdX/loJWb7TcXFqONvb29tH+AxZSrbmK11eoQP55xGHuM7tqV3MYdn9GQAXmyPJCV4IhxVlDN77F53EBJ7L3PH+bKukFw5oiNLJFP90XzS76iXhpWbsaCG2gVx5w4R5FnXj8NR7s+Xlr1Wa763gsmW4yz2wUKMpeWHfI8OMZUx1pvbmlWWRi61wJPkBrwsM2zUWPBBfokdDTZd+fT/XjCCqhj3GpbeSwN3F5ZfIHFSQc15xX3TCPzt+l2F3jG3+ku5/DdAL6ryOIkbeJuPAkq9ulPfrr2ta99rQWS0yZREUaK9p2In5TmfUQgJRUJFAncpRIogOwunZjSrSKBIoEigSKBIoG7QAKoHYGq1PPS048/Vv+f/sf/Yelg/dZ5Yvc8vbu1+XhtMjmOcoBqMNrE7eba4sry9U996Mm97kJntj/557X/+Q/+aPrnX//68McvX+0TXmgfe4gddITdocYE1Im66DDV75qcZoamqvhulI27QEClC0UC95gEfOHi7QLANHh3tRxrAyYMRHYAVAAGgAV0q5xO27yZuJkZ3bw25t4BbnnbAKsFVk8U+1hekIYr4BxcASUEJlwPECLkmUxwGxwP0wgXw//7L76ePvJv/lVqD3qpD5hyVUPBhu+7ZQxsn8tmyy+vC0QC1LC3boHZFMsqjwU2tqH1ka6SJsGI9Xi/AZ3SHa/qT/7c8IGhDusmY8CWsF7jPBYXMKi/XyJglFZw2KRhFztOrS5qky6EWKARzJ1x8dGizSagBVQF3NLGTaFw5reN8VTkyvY9DZdN+hcQirIBeqio3cR1klU0W/wmQlkq03qtDXTqUy5brwn5BEimXF+2yHL81TXcA/O4/LLSYJafX1k6NE/Cx0nQpNt5hHbh8hr9NHf8/qIqMq+TU8ZwNFfWCvxsAgMFeMPBKOYi3wfIMU5EEpZqVb9C5MxLVYeWZTF/c9DJLebP8RBvTfdUIaYunjZN35xbZeDcunnN86YVz++bp5KPcjR5LR/Xw12Vc7rADNVrLfJ2eaaMszeDE/O4jLBso8fN1iLQb5X769zfB35O+v1++9SpU82b6zfxxjzql0E5bea2kD0rqUigSOCelED+ot6TXS+dLhIoEigSKBIoEigSeL8koKKHToECZAvZ8uGHL71c//++/hedR44fP4FLzEME6nl8uL9/BgVmZTTo81t4dY7JqNlpz/YOdlp9lNDnf+Gjo9/59S9uv/raxeuvvXbxpeF49P3f/5M/+9sXrm1vGcfZ6lGXKEns7KxghJKBOom24Z93l1SI7kxzheXOS+W4SOCDLoF4SXxXBDRYObk44iK8BBAWLtLbACNWs5wRsL+hlx/rWwqhJuoLXfIeNJrTfQDLHqBbcNDSjZG9QE3oAf/hjbUgm6kB+IBIUC1WU5x/7VvfTP/17/3z1MYVT6AV76lUhCToEGQYOMo/cUx9fgmmNI5fXMQAsx7svMIay3ICFusx/7wfud55nUKYqJHyM+AWFVJfBmNCLaxfgSe9DFAYr/BNcKaFEgQQ8IUbJ66RzTxWwE2GR5ge8ZEEZFFh5PFYl0GuE8yKPgi5BEUANMYaVmnEGwtoRN1AxoQXIr+C4PtqIHrG7RiEfUPKG6dNsGTfqyTXqoCY12zLMVebn1DrcHw55fPqQ2obQju65RBjruYZqYN+c6Islbl1VmDLAjFX82q1hMufa5Y+PThI+/uH3K/RdyztSAGvyBOrlNrY/Jp1uAVEVKbMncaLATdpT4uxCWaKZIn27atuqtkMj3I8iXcCstFQWJmt2Gwj+hh7QaLwbJ6fvgkxjYOWs/EvFZAXK7IWoAvryboGZDMYGQy4oRNunSkhFFmzy/h6nSbLLTQaI0Dg9Kmnnqpfv3U95n11dbUONKsdDvq3J8kW3i7N5fd2t8v1IoEigZ+/BDJW//n3o/SgSKBIoEigSKBIoEjgLpIAekmkuRo0P0uziy/+uP7hZ546ffn115/BNekj6NKPjUeDh2ez8ePE13kGDeUpLBGeIpj04+1O+/HFXvep2XD40dWF3iPPPPnYuU/8wkdPfuH5Xzk1HQ+WL7z8OpotbknoWDRgsJ2p7aK+GRQ8folXNfxuRKNCZ6qUpHdTpuQpEvigSID3wxfETfyQVo8d4/XsnccVEbhd2+d2B6DzMPvT5PH9WwQiHBOOQAo2m81Wnxq0OFsGgHR4z6QKATK0eiLvUWwnygYkEdYINNy4kgb7++nXvvTFtNzDxRBLLTIBRWQLdIu9QfDNZ7lwkcRtL4Lqzy2+tO5xy0H+M/xpA5R6vQXAE2oNIMRhClh05NP6KhIUsAJLsTolIMY2dOXrdNoR/J4xYjnUCnjXpJ62Qd/J13FPfXX61wQicQbsA5pRvsW5we4FXcKgsDwjX9sVLOlBHSAjT3ORAEGaG955YS7rbwWgZgH+atzHlAkrrEPcPAnnCMjCDzBikum+qvWY4+qxWmNnoYdLYpfA/3AdruVx5L1j9fvnNfe3v4XIhXvzyWfcykUheSWqifptQ+Fp2WcdlZXWkRwtFdAqu0la6xD30NcvXko31zfTzt5hurm5jd88AFQS6LODjIIeWfc82U7AMazvdHXk2Yq5Eo4BmwImVpDPPtgXk1ZuGb7ZZ+aIsm6tdnazFNB63zEwujzmaIs2nCf6wk0MCEdCXeOPWTdQuHaR/RY9bHOtibPlARl1q+TRnhxubWxsXr9+fcRCBBOh2NIy61lA055//vnahQsXaoBimyupSKBI4D6QQAFk98EkliEUCRQJFAkUCRQJvNcS8H/7d/yPX0MKVZTp1t7+4OBgr7W80H2k3ah9dG935+l2s3G+1+30jh1brZ08fiItLHRRcHRhmhJEuZMWlhZZGK+5zC/hT4xHgLRa+uSnn/3Yc7/76194/KMPn0tbN6/dXN85YHWwMG6gZQPzsMgbaiL7HN+ag5+UVHaqdOdxda3siwQ+qBLwfQCW+IK4sUpfK505c2aZl/oUd3i/m4fNRmsJy6fHuH82IMF0uoTV0yq+ZEOAynXeZ4JC1U9ihnMKCOE3gfiB4oaptqMBxwRlpttgJk7DLbKGiyTx/tPqYjd9+uMfS8P+PgCJDwtZAnroSkee6KuQgzTpEx8M2DEyNhhlB+zNG5Zq3G+3ummR4OmuFqkFlOZZopH4fvFD6zGTnMw+ZSdIYFYDKAZU6XYXAo4JaHSXtKB9osNpMmDlyCFwxnJc84Pk8rxCMzoRUAxaRz7gFUALqpJqnDdGwK0B1l8MwfwCMe8LwGoca67nufVorSaJHB3sp+HhQRqyGuQEQLTPipB9YOKQ+wKo0WgYVmgrKytJICggw6aJgQmaGJXjtH42m3SsHufpRsYex3mWq0P0moqgv5SI+xakT3FMHzmjjPKzHotrkaVsPXcjD5Zumxub6eKVa+nmrfXUxy11fXsXCzj7onWb9ZCXv1rCVd3wuoCs2+6mDitz2l+3fWOZIU+WR+UfHNpzLPPWbF8OFSyKi8ZfE04GYMPllcB5xLQbEyjP2HI0OJeB7WjJ596HlmeUR0k5yLiQQaNxgAwvcb5FY04HXa8bd29kSD6e+73XL16+sbd/gBfpIK3dulU7c+pk7WB/f/o33/1bO2h9IS7KvnNSbG4lFQkUCdy1EvC7WFKRQJFAkUCRQJFAkUCRwDtJIGuZqAL+335j4+bBf/Nf/sv64GD//NLiwkcWF3orHawZAGQH3U4XfS6UuVG31x3jcjPpdjroNLMGv4nvLC4urmBPcLo+mTzaazYe+9ATTyx86Qu/2kPR6fz4hZfUfQb852SI1xOEjfbUc3DAodnq/yzvShFRmcoK4jsNq9wrErj/JeB7IHyYpzhYXFyq+S5yb4lXDIJDRPSUTvG2Pc01ARmchNhMWJDxUk6wriJIf30MajlBnmNAAz8Fk6nLMKLyc+/IUswGgAvRppZj3tPqy+vaHW3dWkv/5MufTzMWB+QtDchhnDHdKHVlNMaYZaaUEWwIxKwH7MRKicATzwEcXusAWFpt4BawyzICHeHLBOs0V6Q0r9exHQKMUC/tNbAac5VEFuCMfubYYQwH66UGFl9TrNjqY0EY44DQaDFWAa0aeSbE2pqxjYV3ACHLTTmeHPYDjFk+4FofmMcYxofkY2yjg8MAZGP2gr/BHoZLAJ3t9fW0u8G2tZmuXb6arrPIyaWLrwOc1rAg6wOL8hjCekw4xhZxz3RRxHoKIcW3TvkyZyF391XyFxXK2aQraOSZ31QedybPtfwK3OM3VJmSbj8/1E+R6tzxbW3vpFdfv5R2gVu7WJBt7OwYqg38hNQBkfHAUVcFNWOeaEdX0hZgUtDl6p7OlfObn5VsBTeZcydBp21W4wsexfkCdeiiicVy9FWY6IgqS7LcluOuBxANl9eImcnThAVkwLN63RWY16l7j4eeyzylGXiNefYPW63mFs/T7t7e7p6yoJ81/s1rPPPMM7WrV6+Zn9wxSm+/c3qjuN85b7lbJFAk8HORgP/hLKlIoEigSKBIoEigSKBI4J0koFmHwZbr/G5+tjuYDV5+7fWvf/YXf+EYfidPLqwsnz51bLXZbrfqE36Lv7x6rEEcsrqK7mgyjBXD2k3Wfqu3ahN+A+9v/FWgUV7OoK7+Buu/Pftv/8Xvvvpf/NZv/OVff+s7f/i//8ff/5sXLq+r9xHY21+4zyJUD6qoK16icPnnJycVnZKKBD7oErjjPaheiMbK8jIxxSYsINjazzDAqFIzlnasE7Bfi7KAEdCvBuGxiLKf0jIwAXxUO4Rj7GASujAcDrX0jCSIEDaE9Q8ZTEHTeYmFB77v2pYJPF6/sZH+6pvfSV9+7pNAoz5lcCvku4C1DnUAu4jZ5QqTwhAIHOUIjG/vqMfNNiAeOXaVkIh2hSt+MHR79NhYU1MsufxeCEW0ijIQvkHyZwAtDgLMGJLMQPMKhriKAazqwB1W6QSyGXSelRXpm2BsBMyaaslGH7Q8Ggn0vA+o0yLN9pXDCBBXM8A8tTpum6NjXM+upgIgx+ZCAsSvSltbG2ltbS2tb26ky9fX0tYeLorTUVo5tpw+85lPp3OLWLkBgQR6/gaB5kkZ9HlNOQuYQj4APeN7aU0VMlEuyg2Nzzk11pll62Gh9UboZK1KjIJkmd/LjeW5UErysrimNRkzwzd+yHgG/FLEc8dvP3yabMrfagTUomZrhy3Z8wChujzSDBnoHxWPsK4bAk2Fm0LOSp6OI+aUfPbd+pw/05g5ngAzXVzB36YQBzPmPWRBPyLWGfdyXwGfAFUfBuaF9WXsb/SQ3+BMT3NtA/B6i+dpOh5OcC8eHXDtEPkOsLZcZaXO2fr6+gbNjjY3N5vPPfdc6zOf+tTsa9/4Bku9xnOncGN27Ntbpne++5ZFysUigSKBn60Eqt/G/mxbLa0VCRQJFAkUCRQJFAnc9RIIReSNvXSlSdXIycs//sHs3/y3/3qt02rPUHSWsUY5jcXYIgoHYXooSSIuC/pFvYEShf5QR8ecmletZMhv9MNMhF/hL6LXnGnVps90642TH376ie4XPvf8wrGVxe4P/+6FOvregIXdRuh/sjdVM1W90Gro2tuqGzT/xp6XsyKBD6AE5u+BL8PRC4F7XnN1eXURQNbjveR9rB2Qz3fpJDGaHuTaCV6fHqBgBSiklVkL9+ghNQxgC1qaASJqQgXCo1NtjTVtASWc10Z5H3DItgUVATfIF9CCva6WkI30+V95PoMwQFO4uumSB/fQkgxqFVBDiMRHBIsk4AkgZspesGFnjcFlUPgGFmR8RwK8C5DCKkqXR13qADJwq2zlRUD3FuAsYn+Rb4wLpbG/Rn32mDxNDllMAKuvMdBKcKd1GMsWYg0G6NcaTKsx3B91mdQaDdoU8dE0NrJfupcCDcMCasL5gONDLKIwPSKQ/WHa3toOF0KtpNbXb6Wdnd20hfXYtatX0oVXXkmvvvp6unZrP+0cuorlLD3zzJPpwQcfSCurq7hVZldEx9TuYTXHLxnCegwZu2hAJWsF46dP5BQACDjkPSGUe3LHfCgT58MU9+PIY4kVezJYh+fCxbCQ8hpl3CaM3Xkd9A/TjbVb6drNG8wREJHrNze20yHQKgE6EU3AMrvgoyLQMw6YwC/HHsvzZn2CTyBUfl7sB4W0/LJt+5A/99UzhYy4p/UflBf55IUQBKq4BDM1oD7K+FzyPOfni7Z1RxUmAimjRyETeBl7t23yXmZ8uxzze5sa/4DVr7PfQGz1XpfFZ/CzpCyex+Ma75FWZLNXX3sNA0KgbUlFAkUC94UECiC7L6axDKJIoEigSKBIoEjgZyMB1K0JekdtQGyeP/uTP+n/q9/7vddXllaHjU77AeIaPeJqbc12a4wGMSWOS0MFyXhHWo60Oh1+yU9UHitQH0H74LfzePTgjsU1YuucQHF6qtNu/tKHnnj0w7/9lS8sPHp6ZXvrxrX1nZ0+ik2M0Z/qd1YdRipqOm9OWg6oDKLiccuN3CUVCXwwJXD0ivBOpvPnzjWBOl1AAHHo2xNcDgeyBM6XgBdnAVKnAd3HgU3HgQGLiKxGvK4+Ma/wIZwZ4EkzIX3nmkAYTXl0MROI65+WIYpWSLxyghYhhLBDaOFbq6XY3u5WeHIcOQAAIABJREFU+tQnP5FYvINrADLeUT4ZESNKl0ABGYHUA6YYuN33WcssVsEN+OZ7LfjAVdTvTXxj6rhORv1+GGzbTTMm4FeTKg2yP9zdT/1tYnvtAmKAXgfrW5wT92sfEAYgG7OP+GEAnjHujUPOxwC0+NoAXgzSb3yscNlrtaPPWlExUOkP6B6SQn+IbpUGjHUquFtaTK3FxdTAEqyGBVOD+GGrp06nY6dPpTbxGid80W4AzG4Q3F6utLickM0vpF/6pWfT8RMnU6/TC3dEx9si1pYupcKl/N1kXPFh9EMqDLOrGUpymr9/MfvOA9M2B0fir9sJCIWwtHhzRU3b8W5YEXpsfc4rZV2NlDtcE1SO09bOdrpx83o6AJTZj/6AGGSbO2kPGAm1JH/uj23bJr2Ij7erfToG48B5zxhrh8RgM0C/YM6B+NwIR6P7XPNRQ7zxbAR05dlqMgeugIn5MnLpcD9b2VlIWDmmjwJM22kJ56iAemMQgFiGNZsyXn5v0+iyv9GoNV/A4vAWA1ygHAH70y5y3SJbn3+oDhaXFvcODg94lGfTK1evKYra8ZMnEgH8+Scs9/S2XMtRkUCRwL0ogQLI7sVZK30uEigSKBIoEigS+PlIQJ6l7tJChensHg7GP/rBDw5/+7d/6zquRqhYs2ViFR2jawtqHMQvQglqjlBCIig4Snf85T76bt2Y1+qvqD2zYafVQv1kwbh6fQWzkofa9fTUQqu5+rEPfWjx87/6KwurLHv3/e/9aIiuc4gabHBwta0me/4vo1p3W+ULRYXK1F5i5+EdR3FafhQJfAAl0Fvo1Y/hAj0ajuUEvIdBV4YBAGq1VfDFU1x/HEulZfYdAFjP17fVaruMYvgXcr3NNS3IxBVChhn5IN+YZ5EERhwDSPxWZGjguZsQTNgywBrr4YceSB/DSmrcZ8HA8EMU0Gg5ZgArLYCoIqBPLeoUsFnH2Do4jpUcgU26N9ZxaZTGmF+XStcjMLC+JqiCsP7Oftq9tZEGWHIJvLQeG+2zSCF1gZrCddIVKA2aPxPuYAE21p2S8tRCfXxNIlYWe+o3QL7fN+Ns4W4KYGLoiHLWaqYhX8IaQGYGAJoRI6vOCpsNrL6Wj59Mx06dSqfPn09dV6MEdu0f7IUF2euXLiXIS1pebqfPPvdpXCs/lc6dO58WAgAyPuXAxi8iaAb3UupVtk5fBSHjW8cPLfDIGrKyr1UKqOQ3kcH4G4acGDsHQimvI/EAmdgBz+97zXt5Ls1rPUJMXUV3iDe2zwIDA+TJ5bSPddzN9e20DWzUPX5KH3nMoo6AZMgm3GgBW1rDucWcAj73WZRAmVbPTMAxx+hg6IMWcT4Xtm+yHJaNsVcexjQLl9OYrPwcBrx0vNShFZry8lgZCXc5Zppa7OpakK1jfXaB/RZZF2hicS6Xfe5ucr5FG3RxMtvc3GDF5fp0bX2t9tGPfrR26dKlCF6WZWjvSioSKBK4VyVQANm9OnOl30UCRQJFAkUCRQI/BwmoLgme+KuWUru8tj773vf+bu+3fvM3XyX+zw5K0Eksxh7lJrqI7iyNMQcz3GfUckBkKigyLVykWjg8NYn2QzwYNBaVlPrYoNdWXK+3Wp3WGRSej7RbjY9/5JmnHvhnX/3y4XPPfuT1K69dmK7toFSjJ6K/aoVG0BrKVDqd5fmjTYSKVd7YlVQk8AGTQAUb5sNunDt7tgtg4D1sjoQCAIc2sMTVKQ+AA+d4Jz9DmScbLcL+1QgfOBprQdZrtpoAgZpluF3TFLTDm9XAqsilAAVYcGuNtLJrpEH0TZ5rxAUXCfChG6LvoyBBN8PPfvKXsJBqAqwGET8M0pbAFXQnKHq804KRGZ10bxww99YrINP10GFoOeRYPdbFThc+vgrpcGOXAPgbBMAnrheWZCMC5g+0EgPICVc6gDWvt1ltd8zeVRCH5GG5wgBRdkC3UU4Y3TxOFjBnYjvApzEfH53rhEFjrZMAYVqKTWm/1sPya2U1rZ45m0498EDAsaXjx+gb4Azrpu1bN9ONi6+mNVwsb22spXNnTqbnP/uZ9OzHnk2PPflU6i0v4z5KPbSNeR9rjWYopEWuMEi53wZkSjvDrwzFPM6QMb6Gyp8Pph9hP5PeM9UETFxQbgGwyHDndzRnsi7kH/OW59Q8ukTu7O1EYH08D3GBnaQ9ZHdrczfd2j1APjnYv+6zzk1OGXgBXMM1UqBVuaXqhurz4bc7W+iBLgV89F3XSVrmcc2Q1OfH8XsbeBX52gBJFzCwLUGbaYiLrE37b5EHlGDe7ZfPoOMOCznFYrltst6kQYPxew3zxlmH64cIaY1/u7awKuOZn7TW1m+JXuFss9najRu1X/vyr9UuXHjJEHclFQkUCdzjEuBrUVKRQJFAkUCRQJFAkUCRwLuWgLquZhXqFwQUS50rN9fGL3z/e/tf+cpXLvYWuhh6TFG85V+tBdykOig5TfUZFEO1ltBc8FBhIUvDiuGIg2kGx6GpoByNsZBA5wylR7cXrFrSIxhsPNhtNbpPPfJw85eefXbv29/+1sHW3mCIbqRXkj1qosNV/6+JS+96RCVjkcD9K4GKTKSFhYXmiRMnusCsOnxkxHsKhW51gA0DQMWAd834Y58EJpyDaAkJhrg3rpJvhXwSbMqAqmo1XlkcJbUYw7qMfC2uaUFWIy+XQAduHAsmhB6UjfNw8QPGCCu2gFZPPf5wevShBwOKkTEsm7SQ8oXWYszOU3cGHoCWEVZddRa1DTACFOsZgwxg5PfCtiQUYiBBWB9I08el8gAXyj4xxYjKzrAI6k99umwau0qrIq2YRlqUYRElCCJWIigG0EetgimRDXfSAW6ABKAivtYk7bPt0V/WpWTJXcrzgaov40a5spR6J06k5dNn0rGz59LqaV0pT6YWFmMNrMsEP3Ws1q69ciH9P//pD9Llly8A4/rp4QceTB/58IfT008/nU6ePJW6WI5BYMKFUDjXaPlJ5euIDOyvY3VTYP5Rnn70lL2JU47z6pdxKf+I8SrPDM8sk8t6rSo3Lxxyz3mpE3kxs8xhrj+7RB6mPay+BGX7h/uAyykx18bpFqtaru8Sq82FCsju3LuZ3GfLsbxQi2UEni5WoLWXxybzmFdoF/Hp4ncot6GreexbtQnShIZC0xgL7QrVwi10/kxan3Nu3WSyCgfjM1vj+bbcHle1FNsgL7+B4VK9RlT/dIhcr3F/mz0LLtdbkOPhwcH+uAEEdGEB+o8hYSNizZG/pCKBIoF7WALVfyTv4SGUrhcJFAkUCRQJFAkUCfysJaBmEdoFKqdqy6XrN2d/8md/3P+tf/LVV8+cOnlxf2cbpWJ6HAXinBm1UJhgikFcG1f8amLCopkARCsrZiovKKv8ct7YQ2SjANysrjuVVhKNRmsRXf4Rrn5sZXnh5D/7zd/YunHxwtVXL69FP9BrMcuIPoWGZd9KKhL4oEtAxKAMtJx54vEn8AxstIeDQW1scCYuAwa0/BqBd3jRaud5D5/i3SMKVm0PqxndpM/wLq0AY4aAhKNI5KCJMVtY2XC9i8UYbIovgUAJyOF7bOwn4Q312YWAN77LwjPfVEL7Axb206c/9Um+A6w4SPkjbsGxrpbCr7Dg4nNhiu8Iq04KulrcEzhpgBrtGlRf6y5g13CPWGNsB3tAMmKJQXakHYA44l4FDMH6C4sxu2wfBTnCGvtqHyGB6QDws4tl1PbBQdoFYvXJjFNmGmL9NNK18/jxdPzxR9Pyww+k5QfOpRWsxBYBYstnTmM1djq1AGY9QBc0jo7TikMArG3fuJH+6H/539LWlavp5Mrx9MQjj6bHHn4snT//QDp+8mRaPX6CiQEC8n3Mv0KopU6XkG/UYewuLcqMQ+Z93ReVCQLhmAYcCPL1j+MNUdOsYzQJBMMSa35Dt1HvmT+Sc0Ue6Gd8m71qvVabra4yPMRFN+3t7bIQQcChgJmIDKI6SZvEd7u5tY8MIadAMtsMuVJ1p9lmNdEcM87nxDk21pyQLZ6bmCc+5sxRgCza998Gu+2qos5RlYSB3jMZp84yHWK8uXiBZQWsY4CmoDaDw+yS6XjC8i4vTGEdXKKPtdoBPzYQx1Wau8E5Ye8mALJaH1lf5xwLslh4pra8tHy4t7uDt64x01Jte2d7hgXcXIhVD93bP2X+Fre8XVKRQJHAXSeBAsjuuikpHSoSKBIoEigSKBK4JyQw/18/ejH6Bv/9727tHoy/9pd/0ccC4lWiG22jfPVR4A4J/I0OWze+WA89oYVfCkHDatN2s4n+MkLvQFNB2UGhQY/CWYpfxes6yYlGFBh0TLEUa7CYZW2JrA/ihkWMsknj07/8qdnlKxdnr16+OaQzaMFhdMGuZoy0opXcE49R6eT7IQHek6raOFgC1Jw6dap5cHDQBEbMcFUUkGH1gmO0K1nW8FSu1U7zzj3C9SXeR8JH1RaBFuc47wEf9ngPWe1ybugpZcHQh3wRo0y3NYAYWcIiKN5n3+noB3vhmcdeM2kVxIW0y0qOzz/32XRsqUf8r6EvfdyfBgxxBULqtQzZtZgSkAhC8vIc4aYdKxVaF3SdoPoAMcDY1q31tHHrFvHGBsA6+gHu6eBG6aqG1hF/BCe0NgD2SNUHwBTW60wD+roH+NnA5c+PCv51qXV8NR1nRcmzjz+RTj32SHrgQ8+kM088lpbPnw0g1j22ijulwfgXUpstzFoZSzAY4M0Yl8oJVmzbN26m177//bR1+Wp69Oz59BCWY6dPnk4niE22dOxYWgG6NYBh0L9YndNfIrhCp8BOGQialKNxvHRPdFzKUss3pGyWuF/Jm9Oc5nLXM76al5gP0SltCHCo4ihZm1Z2IVfKRnGEpcRkq30t9JBtf3CIPPOKnT5Sulny70C6eguXVspXrq/K2X4GMGMMzkiVhGOuUGqq+ib4cvPcefdxEbjGH67ZpskxuPnc+Fx0u71wndXSLgfozxZqVb7s4k+/kCn16x4cIpvDOK0kD2nvGsjsMmX6tLPAfkZdG1zfURBY0fFLnlqff8fGgDHbtw6H+BapGufb3H6LEuVSkUCRwM9XAgWQ/XzlX1ovEigSKBIoEigSuKskENrCP6BH/rdfFWWuXM029/bSv//jP0v/7v/4j9t7+7svP/XE039bxz0Fq7AFFJiHUFxcxlJlFvUCv0oxGD4rWLSEhQRmLOHWRJWeG6OMFkI9wq2LllCaUFSOcfBop9168hc//Myxwd7G9muvXr2qxq/WTvVd+mXXPH1D+oeO7w2Fy0mRwL0ngdDQj584jmVNs3nY7zeBJ7Pdvf0BL0gNa5u27xRc2pBaJ3kZH+X9OsEwdZlcQfc/y9bh+i7ZNaCCc+MVHUwgNQBixmjynOxUDEBg8yQgmUDFP+Z3875JQEKbuKf100KvnT721JOx4oa8Qogh4BG6CSRMAiHhXJW0UBOIWKdJoNPH3e+A78/ajWvpxtUb6dqVa+nm9ZvpAGhG65GvTWB8LbpESS7H6wYtCQDV5+qINo0hxkoG6dzTT6cnf/mX0pOf+ER66CMfSWeffiodf/ThtMDqk8tnTrEUCUHhdelrY3EGsBnTV6GVYEZXzwbAbkTb+4C6Ee6kGxcvp5svXUiznb308Jlz6eypM2l15ViAsQ6umQsAtgarWtawDmtTb6JeIZPunSPGaxuOV7kF6KGvWoApTeaEe/EtDhn7rVTW4cMeNwSU2jMJHDOsCtlFnDDnh7J+Zq2Ntjx07nIe6+K3DwJFrhunbYBFnVvflT/5dg9Gg8gzggzuAgIv3ljnOy6Ics4oFP3RZRS4ybGWYwbKt6ywy1mung3bnAOraJ/nMcY5YeVM87gdATLGY6e8Zpk21n26WRqXzNEc1WkvqNc/1se7kMEbD1yVhyxU0dTl8hamlpfIesgTfZzrHcrtsG3T5xF5eEzqWFTOxmvMrc9lyM/6PXhDipG94Uo5KRIoEri7JeBXtaQigSKBIoEigSKBIoEigZDAm/97/y7EkmOSoU+F8jStGQusBaw6/OFLr2x/92++c/nkqVOXjp04gdHKaLi0sDyZjifELEoE/56hPqn1EjJbUws0DRW+FoGpRyjIocfVCb6D+Rg3OZ8Nyc9KlsSBaTZXuPIUOtHJZz/64faTTzxc++53v7NNiKJDxqA5gjYX/j8na5DzgfwjxvcuRFCyFAnctRKIR974TAClFgHRu/uHB9M+vmG+X1xfABi4gp/LWupa+RDAQCjAaQ3/wHSafY8sWIMGBHP1Sm/usQ25rxVZl7c3/PmEYXMrMvfyiEjkzQf89Ng8EQeLt39z7Vb6lV/+BLwJdzw7RVY/BxmS4Tntt0BCQxJuuAn1dLGskvWNsNIasqLijjGwbq6ldazI9olB5vkBbpbSclecPNSlz/pob0YdmLKmSbcZ7pFnsA57mFhgj37so+ncE4+nlQfPpRbwqr60SLj2NitU8mFhhUdWNaAssIl+RswygZgQCAsqAy626fOQFR4P6cfB2lravHQ17Vy9llpYqy3yfVtdWg4A2CGo/8LKcurgjtlaXkrNntANSzfkwm8PCMzPLww8pj5dEbX2EsIJErWacq88QUaxR1AhEuchrusbScLoKfb+JkOYxjcXefA1pb7IxzhM8x3X4jR+6Fo50XqLvcHvDarv5vmQD67WX1rvGa9twIqhe4NxurrGiqGuTOrnnYcgvuYcOXem289Irtfz/EzkfthHN68JQk30PMBaADXaimshg2xp5jg6rB7qAg26oJpyXLnchveVmUkXS+rnErLjAaNfWpPZOWBwfY1rr7EfIIZTHHe4vsF+HeNmDOW0vjRuX2O0C5DFAo5s/utXUpFAkcD9IIH8lbofRlLGUCRQJFAkUCRQJFAk8FNL4M3/y1eBeMvk5TtuzbOxqxHMCO1LnYwfG/t76Q//37/c/cM//5NLyyurL5w5cfy1HstSUvYh6u7AzKwItVIlWP0JZZXiTawnjLWTV3BD+VOR45f9ZEZtAqOh0xP1iJXvmqsoRI8/fP7Mh//F7/zT3qc/9uTlCz/6we7G/tDV8/BVCl0PQ5E7OsvFf3R607h/Uj22i6L1k7KV+0UC76kE5s97BlQ8s0PgCiCj2e31uoeHOA3CMgQCvV5vCYsYvOmamD3VF0EGAjFXrmRXWyTPaY6XeN+02vF9kjzoebjGvUMARo98S0EvorUanGSGF/SEmPi4UvsVEGbwHnDZSimKFdKM5nh/BTYDrKxOnzqRnnz0EayXhkb8DzBiXozT4t0Pl0HeoyYAxC+AOIK+Uq9WSc1YCED3SYPIE+swPj422wfg9IE5so9D3AKFY3WstE4/+hAxxFZS49hKap1YTV1WkDymCyWWbEtYiDUBVgl4NRVQAcL6WDr1x8P8PaL/WkaNgEJ+6bQYqztO4FGD46bwiPhco7X1dHjtRjrAmm3CQgEIMS0C6HrEyXJsBu1v00YDKLbE+OvsxwAvgrulkRtQDJ9EVzEJq7Ea/WCuGPJ0HscLNY58Uq3YUWes3siJoonEgZZh1bkozWPCyynAeSZ21SF7pzFgnxZbnlFggptqcCE+qlj+EhfOeGBYjmFFNsYd1rnFR5dnbEzstlG6eO0mz5xYTIu9DLByf4CK1KmLq0H0dXetngu/k9bp/s6Un4P8HXWVY+ONxWIBPATeq8orG8FXRwsy6nDzGbCN7BrMkOmLeSxXgTfa4jGOBSUkZhguNgRkF7muWZxWlMgw3WInJBMkQyrrfeLjjbFiTts7OzzrMLNKhnd2vhwXCRQJ3HMSKIDsnpuy0uEigSKBIoEigSKB90cCoQioEPk/fZUCtrdNb7p1R1YNNcKabMIv9MfTWXtKPOztw9H+X3/rO1duXrty6dlnn90lNlkfJWyBaP0rqFYd3Ckb7U5nQpDnKW6VNF3HS4k7Kk2hZGtJ0Kzj/oM1mdYlKCr1uvpkl+zHiKT0ZKs+PfnEw4+kz33u+a0//dM/3d0fTP3VPt1QLZwZjNyEyvRTpDeN++1qClneIZS3y1euFwm8jxKIV9n6hQhLS0uShzbgAMxRHwCWMVbqdHlWSXUVf96lxgn2y+TvAApWOdaCRsuyJhBBl0otbVzh0hX9rNq8S9kYpyY4GwA5CEY20UWzIh2+yVSVXx5hBMZAAccE4k2gRf9gLz2HO2NPyBHAR0spYIp5eX/xZrMtUgYiAUC8T5XW6jfB/hi0n+8IAAkrIt0yuddstMMtUFh2wGqJBJpK5x5/hFUmz6YegKyDO+XCCeJ/nT4BrFpITQDakA8LHw5A3jTtA4F0bzRAvhZj9suh6IponK4aUIjAiqkD7G/sHabD6zfS2oULaevSlTTZ2gOYTRIrjDA2rGOJgyZca2npRDutxV6AsUTcsWkH+KU1my6gAjggUkAs26A9reaESh47ftt2H/f8QVLGbsqiknfe53Ny+4sDK3vD/Up+1ud3N9fm/JKfscXiKchAl0itsgSWwqywJEP25lFGIwDWIeNd29zF1RK+JByb1xZ9RoaRkKN95G8+pc/RTsz3bUsz+x7gK8YpqJu7ZEbZXId5qrFqKakFmZvtBdSjBfdVHtut6sxziSs/eUlEA8A3mNUqOd9kO4CY4Tk7GzCEAdd9tg+5vk9e3Cwbs2Orx1jJc2/mggXzYVpPSUUCRQL3sAQKILuHJ690vUigSKBIoEigSOC9lIAKRFaM8v/1Q4+igbjKvX9IQu9BBYpthvGBWm4Ewn7p8rXBiy+9ePErX/zSd3Go2uDGOdwrH5y3oRYzwz1GZRyFFPcnlJlQXmzeClFOsQJQn/MCWs20PkVpohyWFvWzjVrz6VMEXPqd3/rK1g/+9ttXbq7vaofhuNBqw8ih0te8+PcGVSlR1v7TpqouFbKQ7VyRq67/tPWX8kUC7ySBeM7mT/viwmI6fuxYTSsrLK4mcLEJCj5GTARdClMuYHO93gYIHGM7wa2TXD+DhddJ3rUFXjjhga+SoGCfzdU1dD3TDbNFPmB07QCujaHaqA5HawETgGThjhkB1jXPqd44Y2hp1QMX1wqUgO8H6cEHzqfHH3qA+F2sXun7zH3jXgUUUmPxJSZvVCMwYfP7YFwrXQjbWPM0iUFl7LIeboosAhKQLK+kyHeDP4KRgDt8kpoAqQZuk64O2ep0U2dhAXfHVYgacArYNcJiDMAfIEcLITfb9H024H9XUMaKmV3v6c55+Uq68f0fprUfv5TGGzv8diDhTtlJPeumXT5crGq5kLrGOKN/LQCZlmJkSI3VhTTBapYgWmkMIBPO+cuB+MwhC0EgBCmAIZLhY8Y2twBzXFpvhYByifn3JsMz++u9sLriq+z3NLutepm62Xk//lBNniauIv8Zc2E5XSnxkQ9rLC3nLK/1mNZZQ2QlgHIxAS3YBly7ub6TtvcPkTXd9vOs5RbtxgNwZ3/iOLfpN7/6VsY3n155XsEsr+nGaRsZnEbHIw/PlpnDmlDLMOOQWU63VPumpTKGkgH6fPasQ4hm/dTLLgAu01uXxI7YD5HDJs/gNc4PeAoWEQwzkzY43+DfHIXYunb9+uTy5SvE7xNKxj9zuVPlZ5FAkcA9K4ECyO7ZqSsdLxIoEigSKBIoEnh/JXCkzdpMpTiFIvau21VjiOA3HDTYep5cW1s/fOmFFza/+KUvvILlicrJCr+7P15vNSMekgoscEwlRQsKWo7Ww3pDbQ4thkJ4NaGkqGSTo08OPZIIplwn2Nnw8ZXeQutLn//i8Nvf+uYh1gysvhcxtNUz9VEy1BF/57ohB+9HUtGsUnXMWKtLZV8k8DOTAMCgdpwVEkkaEE0Jei+vkhAYdF/uMOJN8lg3y7Pke5j7DwIIVnlm27wzPsxSBK3EjD92wF7XZQEbzBonQ6w6eXfdN4ESxiprCCdMPvfUrd1QABgAXAYYQhcgDLfSiBURn//0L/NyYiVFmdjiHdJqyzOuAdQsa31aV2kxplVRE8sr4VXEmJLKRN5MxQVInQaxvjo99q20ADwZA78M6K+7YBM3RiHWIit9Gv+QGIn542Ab/qV+/cb1L+1hAbVEHR3OJ1u7afvSpXT9Ry+mm0Cx7YsXUws3zjZxxk5Q13KPFRUFdoCaBm20gHECuRqxz2pYjI1bfN/Y15d7BPxnKsjDFy0+ZPYgZCX84sMWYuBb16rn1SvJ5ggzJMui8QIwKz63IWPmJcsp7ig7J3EOzbgWgBJwZT1VinY8iTYtzzgFTMjETrif4Rqbg+y7Z+O+EteNtQ8wHEH3tvf76eatDeaWquwsfY/vOW1Fv+YNVs/H/JT+8+13Htmiv7TpfFfPiw25SIAyMa+b+fxnwjw+A8pbSzLr8DkxTzwvNJL/vSA/465cLM3PfeGYZWbU43AIwj+9Ts8vUv+A5/o45wrrJnstzHrsO72FxeHa2hrDMOzlkcUkxyUVCRQJ3KsSKIDsXp250u8igSKBIoEigSKB91kCagkVJMsqlFe8pqKRr+STuPxOP6LIPIOaRLpEYO5v/NXXD3/nn371xeWlxc3+8PBUp9N6FCsENO1QonRtIQRPmwXJGsR4QcHGcgyFtjZG61LRwcyEjqjMoBzV9N1BzQ7Fqk4AoelTK4sL53/3q1+dvPrjH669enVtO/pKZgiB///JnkYcWIt9ej/Tkbzez0ZK3UUCbyMBYo3Vzp8/j6WWVj+sjVhj9QuUfJ5LQn4ZCWyGMVMd78M6DKj1AMr+E1T1AO9TjxcMizCDSRmfKSxsNrl3HUCwA8YQSrHkYupStoUrnkGmmsSlYkGAQegZvsfcy6sFWhnfDr8kgi0tb2gLkNRKt27eTE8/9mg6fZJ4XHEZRETDWkppKeZbqkFcvOO85xljUR+wQ1dNs1RujwROz7HI+Fbgxp3axDJrsdeSTkK+olUX9Y52dtPexkbaY5XJHnBMiGZdWrA1a1imAbt6WK2NiSE2WN9K/Rtrac/VKH/w43Tlu996R1tlAAAgAElEQVRLmz9+MU2vryWWB01L5Ftu9dLC4mJaJAi/MMxxNQwYT38b1K+FWA3rsTEwbNrl3jEXAMDaiRUxtRoD5YTVnGONxKAEPw7ecToWFzDwdkChEFTOWl2Pszn38vvttycs0CgUx84Bf6wkA0vmIuRrBkpzbDnhl99a44qZxoBMU6xmydyNcbXUEst5pGI2Le/GALJp2mRxhOvEYMMnkbqRpSDO9qjb1Si1BOT5of1cH89H3PO+yXOT/XUTZgUAow4hoGWj3XleoZ1FLcfCrGy47gb40r2SeGlzUCvEizYcJ+lNkKxqF6NmrCFrtWvI+Cp7fIZnyzznTFFtjV7t8zh3qV93/z4wbniKZ3Y46NexpssDyNWXn0UCRQL3oAQKILsHJ610uUigSKBIoEigSOBnJQEVJZWoKnnuH5UzdmpY7zaZM8wbOOiy9da3d4ff+fY3+48/8cQrYzVrtJVmA9+l6WwBJZjVxFBAssZEKKBpjVhk6IhZs1FJViHDtUp1Ua1HOjbCfoUF6qZopLXudDJ6mphGC7/25S9OX/zxjw5fv3Jzk9L4SamLojFbLqfQH9/tQEq+IoF7TQJCMd3OiBmFlzKUa0ykKyzIAArGFRMMuFAibpdNY4+d58V+kmtnzMsrSJZZm/yAsAhSfot7Vzjf5T3qcP8Y8li0Po5bmNO0AQWubmlZgUR+ackk5PCa34+AXro6AjIEF7h7pq2NtfTcp345tQEqIJMAVRGEPmrI1QQcmX944jvAN8E71TfJYy3LRrg+TkeAkxHtwXZavO41vkAtMmjO2sDSbIE2GwCdGS6Ee9vbacIqjF0Ay2KzA/oYpPHeftoH5l/6wQvp5quvppsvXUjrr11Mhzdupfr+flqFtS/QnsBNd8oue6FLU8swxwWomQHy60IyV+nUrRIXzhlwrL7UY+XKhTTD+m1IjLWATXNAJDh0nLoDmpBtADI+doyczs+v+W3O8EvwxC8O5tcpwVEGXZW8FVkGRNw9+o4iO+rmVgZHUcrjHHesglBaepnHD7j1CZzsn3NYlZ8ib77ZsSjC2uZOurW1Q/w2fh/CGHheHAR//WZrVkablDWGmck6Yl4BajFW8lvGa577jChXR2XbLCUZ9yxrPcoECQXctBxAOKzIvO8z5wqn5otBWIatqtf83OO0hmVlU9dhBSwNXCPjVfZD7i+bn7TOfidaRUjEuxs9+eSTkx6x5C68cuEI2pmxpCKBIoF7UwLVfwzvzd6XXhcJFAkUCRQJFAkUCbyvElCRMIVqwB4Vs9Ix4pqqqX+qfJH5jh+Wq8recdmLqD5phhI1+19//49H/+e//0+vDkeTS48/8NCg02wRGDydtlLBGMqc8WAAYJqNhTVKNv8ikzGMbN1V+tB40KVx6KFAVhuxqZjNHoQEnPv1L/5qb3vt+taFVy6p8Fg16nGtS990yAqN8y37+YZOl5MigXtTAoIGrMdqCwsLWIP5uItaNMYKAsM7Q6By3iVOF7iGBVl6hHwG5w/fMVzqFuEBrm5pMP+b8ARiM9V0qTzFe+e7qgUZC2tM4E0TLMgmDWKR1WyL/PENiG8BxwKJGk7O8oZOG0hEQH1jCwpObhHL68knnkgPuKojFku6N8o1oh7BEjDLFGDMuqyEVCG4yAdcMxC+gfqbuCTOMOo52DlIjRmWZAy3LaSjHgi8UdlTk/pbbDNgzgggtn3terr60ktsL6fda9fSAZZtTQBaG6u0Rn8YlmKrrETZo65FXPkWDLiv1RKLAgD5U2+hl8cjhALsuLVdFRNoNjPe2EovAFnTPW6WU6bCOF8YyYaslI9gDOCfZcUYAwA5Vr9WDDY+hZzG6LnuuXLywyYuUubzu/O9N3NimuYHfIRpNGbHNqjAcvbFHFqKCb20wFLqOc5ZngstB2Ne+GF/Z1h1uTpkg7EOgFe7uFhqQbZDoH4BmYCLyqOfVm59wrUKtNkhQZbzZ4pnJPqiZRgx3+bB963fPHklVkbKvfx83XbJjLaQgWV0nbWNsCLjWdICT0lglhxt2Bb54zllP6QPh1zSzVIdeYMeX6Ivh/Rihd/OwFRnG5S/xbtwQNsuOFrbB5T+2Z//KR7/+qFWSQs4pXhb7tWdsi8SKBK4uyVQANndPT+ld0UCRQJFAkUCRQJ3hQT8r76p+u9+KFWcqwZU17z/5lSV83pW2iKHap6qbn08q/XQ90YYeQz+7oc/fnXzxo2dT37842OVTZS3FeL1E6AH7ygKw72IjIyehsZinCDrCysUKtD9aK41Y3XG5dpsSNuoNA0C/k8e7DRrxz/zqU+2Tp86Ofrmt76zhl444j9Bxl2y/+rIqm8Uff/THXJ4/xsrLXwgJeAz9ubnjHPjkAkDcKVsqMz7Wuli6Ss15rXBE655gusPsp0EAPCKRDB+rcKOcQ4wg+fgekaJSxwTgyydpex5KupwfQTkGgktsDwyDlnAOJrTPEcgEW6WcczLidta6rJqZCTKjAAxuu0NcFf8/HOfjmD9fj8M8C6yEYzIdlxZUn4hkBGQWZ/3tKAyQD/t8HEhCLtxqAgbNQVuCckoGG94g1BRemfrnI39GMvg4nRpX/jm1Me4FR4c4CNKXvpSIxB9E7DS0NIJOLZicH5gFOZ0gDZiXWnVxPen2+2lNvCrhgUVzqsQFoAQm57fDazGIIEBx1ypsrEIJFvkGnAsIBT91v7JcVSbMvFYWeZrTBb9zd877iEIbnvANUp7DxloOScsq77KlXz8suXs3vMjGrvIq6951Y5763Hhk5Cp7onUz+X4vHrfZHtRRpiHzM3rN5hfcrCK5Sht7+6m68Qg29kHkGGsaynnxg8/v/OIPuvCGRVHjflHVX/mU/MxUc7zsCBj0FqzVZuyqZLHmfcS0g1IKSgLyMhkx5hiXMiKPo8Bf7bVBm66z1AtuVDFmGMtl42tt4v81tizimVYR0647+qtGzzK1UIVDUAcbv9jvHW3GVn0hx9Vx7K8qj6WfZFAkcDdL4ECyO7+OSo9LBIoEigSKBIoErjrJBD/7a90AHo3Vwz+of3MelYuFVW+fOnq5rUrV175zMc/foGI+xh6TB9H1+iiTKvYD7AGq6N843yZLRIsakGVLfS4UJBw7FJNUev3AB0JpbCejrNk30MfevqpB/7lf/47o48/89iLV167MNvY3sdJM7ykVP3usACwgtvKV+5i+VkkcO9KAMW/try8LEDSHxkwMMUNMiy/AAjjIBkEwT/N/fNAZV3Kwu8MGLEM4zrD9QWuGacMODa7iMXMGHChG+Z5wEwXcNDHVXoX9zcMyCZdtpZgwnp4t9j5SmZAI1mPlSeBUq4NKNMxr8zkKoHvP/T4o+mBs2fsI/3lXliS+YJn+VM3L3aOO8Yr7mtOC1gURR0jYEw74JPZhSQtoBiRpMJyLHIzfle37AG8BE9hxUYdbQDXErCrSaOS9g7nHSzruvV2xCLTXpWlPsP1s9frgtcaWCrhVon7qiBvYXE5XCqbWJjVtHYibx04ZuwxGkttVqtsANKMNxaxvPKHij76ocpf0eqYwd++xjgQX3zf4nsWnyZcUEOelAs5CRKZGevUUirqy2BMGXDVSmKvlZlzwVeTc7+bWqBlODbjlw8T44ux8qPesfER9X7klGlZmjnhZ7ZGy3HSvDai7AGAce/gMG1t72BJNggo5gR7P3+ZAYPkqyBc9UxUEMtxsoYEeZlv+hznPCcsLBGgzPYFZOaPvnBuHpNWgx7ZVszLfPEGARtPV8jcBQZC9pRT1ngRs/HvCY1hYaYg4JpNQe8+K74eMtohz0yfevdoaI98xCerH9IQGDXVcBOdnTl7Zry9tTM9PHTtCtN8tPN+5Qe36lnOUX4WCRQJ3J0SKIDs7pyX0qsigSKBIoEigSKBe0oCqnb+yQrYO3ddZYat0hbUglQn2hxo1NF//cq1jRuXXn/lk5/45I4KIG5WpxuspodiiMKt0UptimmYgZH0ekHZydZkLZRQrB1mrtCHUoMxyBj1tDZGAddwgRBHzROdZvPhVm229MwTj02++ptfufb1b3yjf2tzd0hGojSFJZn/N1K7KalI4J6XQAUOHAhQqba0tGQMMt8dAQPxw+A+YdkFfG40sZBpdClznEsueSkQg+6k4wBoLcV0o5QAAMcm16mH27WTnJ/kPTPeGAAh7bKvATCWyGNMMm7H+2TeI0AmlOAMQAGc4B3202FeukXcsHHa3lhPn3v+OWJ68U4DNPxa8I6Ga1zUOV8w0ON5G9zP7tbCjoBNfimouw0sk8T7FRizyqJxyAwaLwzzI6QFmDDF+nXBE6C52qUWTz32xirrUAcdCRfzLsBL6zHzGhCepQvCtbBNHa7YCH1kNUrGoRsf4GzWId/qUmoSjL/BeEYsiaklmCCrSkIix8F3Lqyr3Cs1RhBjIbffzNiEhh67dwBa4t1RVVTpfcFfFj3ZzM+Ze5MWaPkg1+lH2D5laAVAAkApdy6Rl75RLurk2GRf7bMB803e8zsMIGUly1G6tbmNFdlBIs5kBO0XHsYikMjMvPPnL8re+cN6ve/wrd9nxGvKWSsvr5lw3w1I5j2T9YUM/dKTtB60ng5zFXCMGG/mJdSl74EdPhqD962GPY89f4HAyGdAewfUq3v/IRl2qXYHsMZ70jAmWWzkQWQTDAYbNV06b1y/QbZ5p+zIUapmKPfv6HI5KBIoErjrJFAA2V03JaVDRQJFAkUCRQJFAveeBOK//So2HPAzlLG3GsWb1QSVGJI/PLSaUHFeu3rDwPrXn//UZ14k0P4BLiwPzWaTk2gjliAGOL/UR42ygIXrKLKqJShUanJhzVFvElmI0whejeajAsg6cAQhbxJjqfZ0u93q/Ge/9dVX/u5vv71P/H4V1q6qE3/ycm3UW1KRwL0ogfl79eauC8dCkUenhyc0dIsUgOEKGQp/H8gkEFjl2iNsp3mfDMK/Agg5y2slPHMFy6sUFoThadjA0oxVLMOHrzbg/YeTTDu4/a1gWQMg853MlmjsA5Cx46LxtVRDADnECxN+mLA9i/06K0uePXcm/eJHPwzUOiTGIGCLP7pW1/H8FHxRG++8dkwAci3ISHXAlaskCkwCvHGHhgJ2aV2G7RygbJpGQJxAYbz0fAfiwxMWZViP0TOsy7AaE35Bzdt8WyArWCc1sxum9AaiZDwsoYwwxlUU9dvUggqvTklbqmMp1lpdTK2VReKO4UqKe+XYviGUsI7Kwol+h40d58I66/QrKJhSVo7QscanSdFxTdgT46dZkA6j9EtIon6hmLHV3B+lXDzXY53Ur2tm5Jr3Q+hkzLGICwZIijbjc0qfkIdJBOn3VhlX/QhZU6egaQ/rsYPDQQCyDSzItnb204gxGV8tvtHk80MrTBNUVWDLuj2uUp5PW8rJurus/mlSPiMMHoVzI1YZ9TxGMpeNHRTAupKlv2Bp4wbrsyBIVG5ugkCfh6o+Qa0ja+Iei9UY3//akHr75B2wP6S/e/zToltln21A264uMOB4hOsnIdhmrdXV5dYjjzyS1tc3MMDz9p3pTfNx561yXCRQJHBXSaAAsrtqOkpnigSKBIoEigSKBO5tCWT1iTGoCL1FuvOqig3JS7pyhQGDKguBXLpsjZtrG/3XX3p57Vd+5bOXqa45m47PovAcR8PBywnNzawo3/z2vs4KlyhhWal0NTgUZc+oheX5xoaOCQVomFWixgI68ENYuZxttxrjzz3//I2//utv7Nza3ItIRXM1TY2d6u/sMVdKKhK4ByUwf45rQIna4uIiDzYB9adTPAnnL2FNu6o0YBVZyRmLZMyeYG8cMl9S6E7tDC9Uj3qEBEIyg5kDJ7B1IvEKa0Hmu9aijUXiiWlB5ksYyfbZ7gBk8+vsBDFCHt3mxsSwEh6NATTXCZD/pc99Ni0BmoQ3BuwXnGi5JfQWqPh6BiCKOrDcMo8wKayrBEnUT35hCt8JwBHXdLUUjsyBifBE67MW7nhabhlwP+Jl0YdGWKXFJyognithhsVW/rTYeQAf5QEyI9oAyqca9UDXAo6lBQL4r/awGsN6LdPD6HsePd10/PbRCyEs6suyirqVm23M5RfFkHOcZ7FzbOkYi18u4ZhFcj3Wb7IakyDI8lEHMq/u+81UdhmOZYhnvX5mhVPCOttzT+moy/zW4zwIorw65nh3fy9t7+ymbQL1b2FFNkVmzhziJI/jCWvGmG8rijHesfea9dque9t1E6JWINWafF6szH3+5yCqPsqfoRqWgZSt5Gd9bvGsRfkM3JSLdQPV/LdIk8VYzZKyPteubtlnnLhW1oRmQjJAchKijTn3nWkOB6P6+QfOTU6ePDm5cOFlhzGXuoclFQkUCdwrEiiA7F6ZqdLPIoEigSKBIoEigfdQAuIllaZqs2r/N19t/9imVJIqpesn1YFeoYFXpKoMikfYoqBLaXQwu3TrVvrRCz/c/Pxnn3u9TdyX0WSE9df0LLfUfl1hz1Gg96LIoeBg0SJt85La+FxZwgIErZbm7Fvo09F2vX6a8k8eW11e/fUvfX7j+9/7ztWra9tVfwRkdkut8+3TTyuwt6+53CkSeM8l4HPfbrdZ6II1HbEmE3Kg3EuahAISkUXcyB7g3XqAUxbICBizRDneubRoFtIO+03KAQx41QjnxbmWaB1esx4gQUDWo27CeGVo44vO+2ioLPILsDLYwTMN32fUETkcr3RYNgm7ybe9uRmB8j/+7LPck98BxXC/tKwQiU9EWDZFE5xFwpJLGIYJqZCcjwP1ksRuAp+oAyup0QCXO861FNOSTbguZNfyyGwClxyOiiK05UdD4NKk78qg0XQ8WCrhpmndwrf4mGGNVmO1ytoiVku6VC53WfqAW1gmjViVM6y2aCsS36dqVU6/MkKasNAS6NCP+GDZPH8sgbzjY1SNJOqYyyJGiSBU7OZzFOUtYxJqed2+IubYHJfzr8yNyeVxBcj4CocMiFfPuBkAeV1pVJqXLc+4j0N8rILJvWZbiz6oKbHHDvuDtKn12PZexCA7HAE8DV8vqGQgjsv2jAlWlb+zzx5Xm/03fwXHvB6QjEEIU7U4tP9kCjk5VvMIQIV2zC6Lh2J5Rt8sF20zToFg5LMc+R2Tc45RMY9pw9hiYyzDDNbvyq26XR6y7dKfsBzjupZlfZ4JhuIoMMnkdTIe2crKyuz82bOza9evh0xtu6QigSKBe0cCfkdLKhIoEigSKBIoEigS+IBJAJ3gDenN52+4+T6dqJjYDdtWAfR8bp0QWjU/Qum+vr4xevXFF7e++PlfvRxWJNPZSXSdU7hmtXH90axh3ETpB4HhxZMDOavwWrF/UFxUgFDOp1oDAOBmRp9W0Wmj+pxCqXlssdNu/PqXvzz+5l99Y7xmTLJ6Gqh2kcf/KwnLTJ6XVCRwT0tA0LO0tAxYACIQjwxF//9n782fJLuuO7+Xe9ZeXd3VK3oDGvtCgKAIStxJUBRFLY4ZSjMehWdxOMIRnrA9vzlsRdj+xT/435G8hK1xBC2JmrFClChxF0A00Oi9q2vNqtwz/fmcm6+6AQIiKGKV7q16+d6767nnLlXnm+ecCzaEkybxnmptmbh1NKiOsB4xocRvebXKyZYVgOlinjRP97vN9TrrSI2aFa5Vrpr1scbmgU3UHmuj9ZVwGz29k0GmBWhB++al3vAFZpKHbKS4pDVEe5F+9cqrhQDZieNrmFeyZGeABis6qgyNJtc6AXosxVPa3HwHIo99wLakQBAEEzpyCGrhD2wGCqkpJggm1iLYpa8qwT1B9zDP4zk0u6hdVdcaeVOdgFbUO0Ztq9KirTnBMUwrMausLwOOufewRfU5DVIQ5jBQ3iAoZv9jn4JGNeMM9kggy/7ZnchDPts2pNJmSu+aRton67H0jN1mjWDf/OIgeGR7XAJigpUBjAHxDPv9GAdr0CF+CQqCpsY7mYMnMc60OwbwE7EL2iDTuvv4ePOEyD00x7Y4yRKt3KIPQCZgyYgFDRKkcbx9KVkiLw3WYSj7m3iceO281c+XQFeiGRNLAFPLBChKOfP77t2rpcks5q6AwlGndRsvQBfl4IH9se641CZEaazeaKid7NxvE6+WmKBwF80zCYWVtS5/eg4GHNsJPVQ3JU/MyToampUHL16Y/OCHP5j0ej06E4Ni0zlkDmQOfAQ4kAGyj8AgZRIzBzIHMgcyBzIH3gsOIO+8Ibz5/Q2JP+eLAs7fFQ5TQ+h6Y877yqrHoDJJcW3j7vT7P/j+7ouf/cJPGjhQRiQ6i+x7MqSPag1AC1FSl/1oOyiIKtga1CQImYt2wo8O8hd5wdnQbkHOUTxF/FtCgeXSfGv+wq9+8fNzL33/u5tXbt69o1jDr8V1fqPklqRXK/45g/097PPPWTZnzxz4+3DgvnX0huICAosLi6wW4eWGOIGKRV4uozbxyxTwmgMcWCT/cYCbU6ywOdIE1F6l0E+4Cy6cJw+mmBM0bIoD1tR8v99fYX01qbIyHs2ALNYPdUPSPZDGhgVihHU0eWMpBgil5pYAt4utP+gXV668Vnzqk8/hwkvwIwEb5i8BK80hBTykR1BJMEZtJesz+In/wihbQ5MrQCbq0h+YdbhfaDbpXmHbbAgBpkQdADk6q3fvsH61qABPIr9moLYh8DRugIJgTlnzlMplTsHkGgOO6axfMIcKyJt2myALosJ4Vdqk0Xp8Io9tpTwJyIpxnGnYmSe9cye7m1P0Utp5MM4dDbSGetgD6ZthSB/MIK+j/7bPzwiASfPVAXyOeqWFfAJzlq9jbhoaZFZC3WpeOX/iNW5q6yVAKuJpbwBItrW9U+xiYrm5vV/0KTMQAGXDtkjq60xjTWAPWso2nBNlCH6T6N3gXWf9aHZFHc4B5lrQU9KEgznoliNoj/E3wPF0vAS/1HJzgkQbtiOPvJHbOOtXYy605iyb2h1BrydX7nH3uU5bhPEBZQ6oF1NM3KyhzRzVTVBYazaqf/Tv/2iwsbGRGEWXKe+VQ+ZA5sBHgAMZIPsIDFImMXMgcyBzIHMgc+Dd5sD9/62HMPZuN/B31KeApOaEIYTCt8+rQodXHUmjffvu1vDlH/+486UvfenKaDzQ6f7xWq1xDIESYTyqDLNMpCfhshCiFJwVoJWHFDwVnOi7yhE4JudIzGlVU5kGjcyPBsNLc43G6he/+HlMn0aDv/7ej7agcthEfqe4oqaom6zjNQVf7udlGf/m+zvJ8+Yy+T1z4L3gAPO+0my2qgINAAbI9q4O1g/CP1eD9bDIu476l2bXUcCjdcAxzM0Ap6dTfAJWbnF5AuYZ8nCv3eV9DzBIE8tV8rQAlqozfCbWC+msTB4BVGyRN4reC75TNiIEYsJsEQf5N29eL1DwLJ58/DHgckAtc6iU5u4RpPNOWZ91BG84rJt2QhMr2kygmyCZNLTwbaazeCscAeTV8R3WG/ZjT2Jj4GCAIYAY2krk0bdWoIh0SG0w6Rvitm1IF+qLraK6OFc0jywCkKGxhGnlmCZ01h8bGHtdWH1yV+E1xQl0QQY/AjEyKAA/8ki7IFfwyX6Z5r7lc6TRJ+ixrIEo3tUG48XKCX5GPfAkIZ/WR/yMXwKN8hqfcelOf0yzjPSocSWopEZuNEOa6f6ESWO0kFqyjMH6vDR71Fn/NidYbu9icglvUeNKdFCZIJ3aZ9ZXjndqJKoJGnwKUGv2RYfPthM0SReXwCPav1FH2S97bj5pLPti3jaafVEndBgsG/2RB05SaDGYl/5XAOJcD0aNiBtCJ39upjqz7BMnYKb2pGtBYExtsoFZSKeBSrF6ZHX06quX1cqUDoOPOWQOZA58BDiQAbKPwCBlEjMHMgcyBzIHMgfeSw4oGpTXe9mOdb9ZTEhiyc9sFXE1iX5qkn3v+9/rfO6zn3kZdYQewutZhI+TwF1qPgwnKIWln2TGFeY4CEENBK0Q7NQgCGEzTHAQaOoVhF2qUDxFCJ1W9Et25guf+eX1//xf/E7v8QtnL7/00o8nW3tdNT6SlAUt9sOrpL98P+zJT0UgoL6hxGHO/JA58H5zAPzYUwHbqs1gTYghYGXaYvI3AM6UDZZZEJxgqelkFT9kFd+Pcml+6SmXG+TZAQxog3xgillMcZy/wTrqATwsjSbjI5wSiA+yiSB0ABWUCeDBNWDblA0wIsz+qExAm4yxntRwqrJeS5BboOzV114tzp8/X5xaPwZkMQxgp9VoBRgTCBjFbUutp3tgiZuGcAw/IOLuBZ5eKC1hZokWWQVzSxyL0V4NTSe0kVi3QGYAZYMAdHoAMEO0n0BIVBMqumg8jdBS4vzOYjqHhtXqQlFdaRdz68tFBWCsQhzO3UJTyhMthbbcIzwEIJY/dKJKZ1e5TPOy3w4F9JAWGckQIBlx8kuwTOhQ2t3H/HH3CWCMJyIpm9owBTgp/JthWG4qPEkgUJSiH5okChINB5h+okVGj6J9eRTmiAJFXPLSNqXdsofAkvURKmhrAZwmnsMn84jR7e93Acn6xa27u3HnMND4lsGKTIdcKuSbB800CTaRNL94IAQviLz/LnjlKZ8eotDA15u0hEknfNZ3Wowr40+pwzp8YJ7TIGrA+CJLX5LQj1l+KT7sI3l9pv+wHq7THsGTX1WzFHndp80b3O8Q5+ASPe2RdY9nT7QcoRFp3HRpebHY3NwqDg72SQq2eM8hcyBz4CPAgVj5HwE6M4mZA5kDmQOZA5kDmQP/ADiQxB/FpNlTGfGmvoVQdi+ulLvUJJu7vrE5/PH3v7//4osvvo5pVA33L+uYxRxFomkq6CK7gXihvBKHi2GWo6CjGgm12G4IngpoSFJoUOiIGTm9MgjBfFrFgrM4Ph2Oz1RH4/Zzzzw7+p1v/O6dP/zf/rDb6XTVJFO+k+o3/A/1U9142wi7kkPmwAfLAcCr6fw87sIAaRDwmwAorQRGVBX8VwEAzrEmjjPVAciKJaCb48ABRwBw1KK5DS0XVsMAACAASURBVBh1izvAmgddoHlWTHeY2WBk43UAtxMAEHMuKy5RBPEGAQxDABneBX7UzprlCYaUgFq5SurVRoBc/WGvuH7tavGZFz7JegZco7wgUcDaAjQ+c6fyAN7i1MtDcMe1b44E8JgPysSuAhhrtTGNxLF+ewm/Ydxbnjy5QLcb7B3zczjdbxRNHe6jhTS/slg0MZ9sYko5f3S1mFtbiufKvM75AdvYa4a4c5OJbhNuFhAJbTzTpn0N0G62P/AacZAdtM9ugE76zNIk0Y0qkuyaT35QRpPKtIvahCBbgGTcbANuA0jpWyuBVwGQQUO0Dzoln9GYTaatEkGagJAAmfwJ80TujlMZLGMw7tDnFwCZnGW/THX7TLa9vd1ir4Mfst0DTrPsFmyu9B/TWbTJAiCTRuoPP2ZWynvMjRm4JZ0lLcb77qU/OAE8TSflhT6+POgg+hfVlIBeKmOfLD8HSBbPtGm75Tzz7rvmmgJuPttOE19nNoCWJVFhhyxgtsnzVa4d8vpliVpmHerY5XlEfAxFoh21M0xX79y5HUCalRFk5j2GRlT+yBzIHPiwceAN/9x92IjL9GQOZA5kDmQOZA5kDvzD5EAS7ZQwFHSUK5Ac7hPG3kaUUKwNKe363a3pt//yLzovfumLryACqUl2Bj82+ElCVkcBRFUDZb5Z1VSXBHOFU4N+h5r1JiY6mFHFIZhI/oAGKIfUdBiOZ+0FFGtOjnrTc+ibtP7Nf/av7vzZt/50+8bGXYvXqUVpKMnBxvzMYLup7Z+ZNWfIHHiPOeAy0MRSp2PMS9EAbc/w5ac/v+oaYMDDCPpnWJMBkLF8TlJE00nzvU68Psg49GJykfKrpHn8q779zgI6nwFAqQE6sNwCsOBQRlYjIdY4j2r5mMbDYXD517FQU8tnjH8wfUF5wqUL2bx3WXv7OH5/8OJFtIEgA6QlNK5IixMrBZQwso695b56owHyBMDDqrUdQR3ID001NbqagF/VVrOYw7l+Q3NJQLKlYyvF0vpKMXdkoVg+fqRY4hIYa6A11lxBcwxn/BXKTTHZrLbQHLOL7FDuMVJxCNq4axkjmITdZTKTdD+SH+WlSEZc1EE+h4VE2Zb2xQQQmd+6Yteknegr7zSW4rTljBxxMzrAQCmy//LRS59jA/x3RaANfXvJD0EkgSnrjbpntAN/sfE6XrXQ+grNK2jxsALri42Z+u27Y9Cj7v3eoNjgNMudThdVX9oF3DItQMPY9yU7gW7SYbvxTmWCp/a7pEnafbd+tcek13dBviGHN0iDeegCOzO/lDdOEFETe3frBnOmgc87EmZ5EwBoPi+DIFn0n345/5qRn4RKxROTNSO+RZ4+bbWhTcxzBz51QIAFg2l56umwfB0zrayuLE9fevllfJTFoElverChHDIHMgc+tBzIANmHdmgyYZkDmQOZA5kDmQP/cDkQwtebuvcG+eGtRQmkGFyPYcSEKVR7Y2t3+IPvfbfzhc9/7gqCGrZioxPcT3BqmV60a8hek6ankakmg7inloACoEJXVI8QpDxFCOFmMpzUxlgckW00Hk5ro8F0EWuui739wdFGrVH9xj/9Rueb/883Oxs7m33KI+oiBoEzWD5qyR+ZAx8ZDqgFNKnMzelGrNpg7akNgxPy6oT34zxfoisnWS+CZwsI/yeI98TKCuU2uL1GPLhX9SxpS7zvc28EQDYe66Rf0CHQD8uQj1UoIJWAi8BawAsEPEgmbwJvNINzbxDYIIH42eJiCVvHazjsX1ldLh48fw40boA2kT6yzKczfTWAkhP+OqZ2gBURb/2B4Lh7hKmjK9e1O9uFLG8e9oY4dZJNoTXfLqpojulLrCL4hTnmRJwFDTNQPOIprdN3ylTok1uMTv+jH7HbEI+Wk/hjDTPO8HtmXwAAuUny7EogEBzinUip4p4ud6fynUffZvziIfhhZSWP6K3ZD0GrVMIoNcYSL3TeP8EkcYTpaNmOfPVSMyvAoaCD0uyPBtuU5hRm7fIivz390z7r61HzVX2jCW520Ro76PWLg/6o2MBhfw/dWy1O+Q6CutK4qoUm7dInLbYT84Rnx8m4krYyvdy/pdO0MRt20CeNVgYfo04/7guCY+YXILMO81qnoJqhrMNn4/kw3xSNNStiGKtqGas5dpd69D1W5xqzAHTe3x0Mh85x/46IUGJlPJqsrCwXnf1OdXdXBbP7WOhbDpkDmQMfWg6wo+eQOZA5kDmQOZA5kDmQOfD+ckCpI10KgUkwvJ8ChZSZ+JoEllmiYu2swMQsN+9uT7/73b/ufOrjz/6kAsI16PceQ1BbNR/CS9/T6agI5TJ9GqEpEcLRPaFIUVkhqQKMNgHyGg+m073d/WLYn1b3Oz0EMKSqSX29dzC8gFLa0m/+2te3X/vbl65fv3mtVH0IdQtaKd/v78ZPPdvTJHb+VFKOyBx4HzkgoDAp5ucXKoANWCyq5OVqECyrCoadQ9hf43nmtL+6DqaAT7Ig8YAym5TRqf8RYlTLGQIezANCn6Rc25MfecbHXxwpSLYEdgiIkT5b+wmksEbTjdeETgDDtepKF2ASfBFcU6NH5/g/efml4tzpk8VRgDJ9STX0IwbUbf6o27LQKRBjOZ2wg1zEwkt7inUCyxAlEKPGqAAVmQFRRMFY8qS5oAXOdFRvfcaHlhj11wHyPHlRuoF5yAtAZxsEaa+hnWo/pFnNMesueZC0mhIlMD32A4pwjz0LmlL+6IHPEbxThnpsRg4aE6dvRkQaz9jP6G8ZJvj4wslcAJF+QeBuG+anZKnQyaAVOpM2IXwMNvhB/71sg+twfMjrfhl8pl3bC1BQoAnASyBOAG6AX7PQIuv2MLHcxw8ZJ2VSobyOOi0rnykXviHtD331SiHNF98CtJMGLxhlHk8/jfLUU84p54Z55J/0GTyiwKGd0nariY844so2AuAjJvKblzLqH0ufY0dOifKwCM3w+aw57+/yvNtotHBLN+VEh8kBdHCqMmAZ/vmok78g0wH+4FBuG1RPrJ9o3bxxs8azji4TUbOu0EAOmQOZAx9CDmSA7EM4KJmkzIHMgcyBzIHMgX88HFBkMZSyQxJgFFbeKsxym6oM6/8xc3c2d4bXLr+0//xzz21w+OTiqN97ADWwpelkVEc40tGR0j/ZNVxClEGQq+ubh3tNky4EtTE+dJTxBr1BZXenW+0eDIq93d5g1J+MDg4GLVRIjh10uifQJxi++MUvH6wsrQy+/Vd/oWA0hAhKolkDUAB9gQi8Fe3Glb19u/QcnznwfnJgYWHR+Y/sTgAKou1FntAgK05wRzOsqi8xTC6rJ1g/nmopYOEpfh3Sza/2mACZ2jPzgAargB5NwQfXML8kgwwIUlGpAEcZfDektT4DSFghAiKaQANXxa4gOKV2kkCPINQY305Xr1wpHn74UrGyuAToAkiGeSRIR+SPdkKzCY0lFHpoNbS5whwwVqogi1BRpAAEUU5aKC/QFVpt+rjynWhBMYGz8JfGs5ph5eUuFf2kLv1iNVtqKLmnJA0oNphIT+0JvLAhUYflEp3SkgAd96EyTlTHen1/cyj5ldqmQ+QTaOJBRiV6jBO6CwBK7S56xo459NRHn/EFZnseViC/BYSCbnavoEdQKdqXT4nWeAjKY1yjTWxq4Zc8pk7qHQ1GmDziz4u4Afe9fX2Q9YrNvR7x1BB8pHyq7F5/ZzHSZICbQZ/glbTZv+AF7z4LkPle5vc0ywhMFkE4x0L6gzbyaZJpKLXkLCcoKM2GAFTJ798E/7BIgeV12O8LedUQYxqO+9CzS5K29ttE0E0QwXSipQ77maLTMTzlmM7KhPGunTx5snL51cs2JEjGLYfMgcyBDzMHMkD2YR6dTFvmQOZA5kDmQObAP3gOhJj3hl6+UyECUUMxF72vYnr1zlbR7+51n7j00M7goFObDPtnO7s7qJhMKv1eF7mwPx2N+nruV/Ir+jh3VlRRsJriF0f5DCWaAMo82e3atdvkGU83N/cAy4bVfg+hb1jMo0m2PBhMVy899HDzd/6Tb+w+ePLM1k9e/nGx2+eUS5QUFIsRc3Xmz69iVrp8ziFz4EPGgcryymrM+zoH9SHcC4YdY/2dAnlYwxfYAvL9MoCEJpdqlc0zxweAD5vM6wP64nF/i5Rps6RQP9Jf2XRxOBw0BDG8BMYIgAsz08oACFwVRM7AAu/lJawjOFYCIC4itcioLOpS20gfZTu7neKVVy4XD164UMyrzaWmFqDKbNmRXXNLYixriIXoTiHwkdqG7lik9Iu4iCSBeqBVgEWgTHDGdE1D1SQTaJE2wSQoJa8aRoAtmCeaN/nyAtChPbXXpmAn9iH1L90lJ0wIpXemVGS65SONchQO0AbORFzQx1Oy4FNbDb5KM3dBsJQe3AMWA4kyPtLJC4AY5ozc1bgzv/yqY55ativgl5T9ojlongGWszEKUumrPHF8HAfrD9BQXpuP916PfZD0EW11+4NigMHhXofTLDf30Cjjhb653aK+Zm9izKxHIMu7PEh8SOCXPIzL+oMW+VSnT+MAu0gNDrmv4/tO2/gEjgWvrJ/xtim/H4HXTc1dKR8grP7QYgyhifrkhXx3vEMbzQjcUmKuO0UDGRw1JpMalQfw9AapG/BjxFzRQb/rAe0xv7Rx3lX05den/pFz5Oknn67euH6j0h/0NGGOvpI/DS4POWQOZA58eDiQAbIPz1hkSjIHMgcyBzIHMgcyB+7jQAgs972/1SOi5FiVLb/nf/jiA+0Lp9ZPN6vFE8N+//HJeLjc6+4DnHUnIGRohm1VJzgVIw0BsRLaFNpH1pB7RmilIBol4RGtsiH+c/rdUVV5prvfn4wHlTFml8jCzWPTMRo20+oiZRvPP/Ns7Ssvvtj9wz/8g+4QtTX+sRIcQyALcY5WPOGvoiObUhiK5LfqS47LHHh/OVCtLi0sgyNVE1pRFCsAB55e+QCzV82wNpPW+zoXJ1tW6wACHYCMXeZ0H0Ff1TPtGzkFc6oz/4XRaDgHMFZL4NghyEK2BHgIpLgAfDcIipRpvgtqpbsLiGcu76NhcsTus+CNWl+7u3vFxs3bxUOXHi7m58TmQOkAfawi8vFeghFhOmk5NKfKYBrrWDiDFSpwZv4EiOlu3YriNEcV6wQ1AJHqAGE+C+4Iv+gAXsClBHas0xDgmH2jjEFTSgNRQVNgLfYF9MYyh+WM4zJdPpUAn7SBElpF0CkgJI/ta9ISA/gCZBJ40nTS/F6hMUY+HSsKAllG3gj2eRcoivbph3fjIszGoXwX5CnrjDjI8T5h38TfFviTQNw4mW/yDDyHI65psbXTCYDs7nanQB+XOPhAXSM1dqUXwDLq8Zngs7wU1Cqffb+fP+Yr4/Q1l3jDxksfpdNyARra71l/OUiVvgIKkr/U7lObL8xOZ2Njnb5bn+NnWU1+adtJKoBMFk5KRpMMEvZp54BL5/0+73FXe0yffY5Kj+c+T3wxM6rcvHGj8sILL1QOuvuVra2tqdprQSdt5ZA5kDnw4eJABsg+XOORqckcyBzIHMgcyBzIHHjnHGggbnmNv/rp54p/9ltfO9+qVf9VZTr5BoLrac1/evjAQVusNux3K739TqXbPcB0civiNUfSRw8SUQiaIZEi2gm4zbXaoU3Was4hNJET+e1gf1hDHqz3u4M2WibLuGc6h6j20NL80tyv/9pXNr7/nb/avbOzFWIsQIDogWJlXRkQMeiehPvO+5dzZg68RxzQp1e92m7NVQECxpiSgUlMjwMgPM77AwA6nnshqrMKIHAEDSpPbh0BofRYHgOEe7VmPAaxzzM+mirLaNWsApIcmleSVgExYAkk08IEfrkSuIQQuOvkneURP+F/DMDmUHuM9AB/WHzqYdUDrEjsUJdHTbJrN24Vt27d5mTLC8Vcu8U6TgCJGkwBUqHKZbszBSKANQty0b4gjsSpTUVkAF2CTJGfugVMKgAqapYGcOZz0MC7YBlX0E9d8CJpjSXy7HLECb5FY7Rk/2w3gtG2zXkiQFbEC4ile8oEBhOqT9bE/mSN8MPi0uyGJG9AmXhTg4t09zLevcZ8EaCWrHugWmPudcJWgnlVeNzggAE13+xXBEElwaXgjTxMdAviBJBDnTwFSd4F/EIbDRNFNbekC3CUdNriTU2zMSjj3i77bXdYbKhBhjrZYDhBqwzTdninFlpZfwBlApVWZA3cHQd5Jggpnc4X49SGMz3GR1oiPWmByaak3ZY06AJocxyZhoKNssexasAD6xOoivZm/Qt/dVbOFf2Wa/KdpqGlwgmaUghuWm/NAEeBMQ+tEDimZkFlrY0nPeJwxTYwb+3uxp3Rt771p5Onnn66/uCDD9YGgIW9nr7+E51BxH0fNuKVQ+ZA5sD7z4HZrvj+N5xbzBzIHMgcyBzIHMgcyBz4RTigGIMY51f2kxc//Yn5px6++HXEqP8Cgeoc8lcFwa2nXIXUxomW44qaDvt7nWJ7e4tT1jrxPEBTTCGyhQ8jtVQ0wVEQNW5+fq7YQQMCI84qppVVLDWVTfGlM66MxpMlhNQzOBC/eNDZPVoZD9pf+fLnKy+99MP6nY2NGgLVAKF8hPiFIzQUJ6iFogYlMv//mr0a9cagYJZD5sC7yYGfnlOVghMsazguZ7nURuFTq1I5C4jwDO/rCPWYjAVIcBoc5igLTY2xPUAZNWZYEfUeQAQn+BX7vLcQ9I8DrC0JXpiO5O/8ruiPSjDFKV1qj5lBWIdYHwOICIDJWIr5bEhVpHTzW4maU4Ik+pmy7mq1Wdy8eaPYurtVPPbYo8UiPtVcpNYR2leUCUf8AF8CYk3MMa33UHPLdPImR/2AcAHQCYQJHiVwLACYmVklMAn10Rd/7BQAh+0IhUf/qDt4zbv30Aab0RLxliGY36AmXDk23svnBAixa8xCyp1Ao9Byov/ydTJF44nninf7xbNAlXnUgBLEKr8EkN2CjwKLAlT2G6qTltvs/bC9kk7KWG9JG4/xbN1hPkp7Pru3hhmngA+bH5hZmFjuH/SLTrdf7HLfwR+ZGmSOg2aaBsu+MaS2gjZoCO086PTu2MS48l7SlDTC0rt9FrQqxzflkUe0Ad3OIcfSvhyOM7QKBjp2QcuM0R4MYVsG6sHMEj1jNMkwpdW/mCbEc64b2tsk3cusc6wPT3LtM74HxI0AIRtqkC0uLI2uXbs6ufL667Unn3yy+q//9b+Z/vEf/zF/QtI4Wfj+UI73/XH5OXMgc+D94UAGyN4fPudWMgcyBzIHMgcyBzIH3j0OqOSlCDrmH5kJRk/rL376k18/f+rENxAaP4ZY2lD+xAG1OlwVhEGkwCTAKiAa9nZ3ix2Bss4eQNleMcZfjmoCbUyo1AypoyigoLm/d4AMXOHb/gFCVXM66GOiibnmaDSo7+3v1CvT8Txy0PFBr/NoZ2fziS99+lOn/8Vvf63+ja9/5eA3vvjZnc+/8PHipR/9KBxV65eIECoI3JNNUUTNkAKes2CUGJI/3xsOzAAYNGFalaXlZdCCaqXeaOA8HP2hSvUhUIBnAFDmAH1uSAGgwCMsnZOsn13KbjA/k9pLteiiULOPWg2Y1WSZjxOATpxeGQCFABlrRPdLaUYLTBgEI7wS0JUACGlCwYd4NYZwnA6eMRG4EKAAeBC4UCPMe4qL6BmgIWBVLa5dv1Xc3dwsnnz80TCjE6RxHUsPFcdlPsEiX6XHS40hoQ0d55fgSwAj8W6emfkk+4b0qallOntPlHHB8hvgi+mG6I9qo7Rn/9X00ocZzIi0aDfIUi9MICbljXJWwWWZ4FWAO5ovzgAoACnTQMLoCxfxgmOCQ4L6pcZY8jUmaJYAKPkmKGR/1J5KtMBjeBTMjy1SWqUlOgHNaZykI8AjCCv7OBlAB4yz/Wgj2oFO+Bt50brzQIXdvf1i70An/V2eu2Fm6TcF6rNJsyH6TQzNUFcCyAJuIq3BaaAB6AWP2NNn88i2A0SE3jaag5qQQnz4DkuVzsA3eUm8WoLWbd9jfOG7/VQ70OA8UCsweEE/wcMi3Q/z+yeEMLW8ypRM8BH93GU67FBxH1dlDGudxTAZkr/HwI9oDyrRXeNPCX0Yd/YPpr2D3uQnr7wS/tNu3rpV6eztWm8OmQOZAx8iDmSA7EM0GJmUzIHMgcyBzIHMgcyBd8QBQSYNo0bKcs88euH8P/8nv/l7rXrlq0hn8wjGfQRkhXPkKcTPmfCHDVEIxS21QZB3Wvgr8tS1XrdbdLl2tjZD48KKVSTT1UwdLRJPNsMchjIohiFBIgSijTZQaEUqQw4a99q1yuhou1l5pBh2T1ZG3eX5enVtbWXh+LNPPnbsE88/v/JH//7/bveH0wHV9iA5/FRzT0erIcuVvbY/OWQOvMccqM7NzeOGSn/jNQT4CopMVU+vfIz7o7Q9Ztm8yr2OjP8U8WdYQ5u8XyV+j0I6JhfDEG2e51oDJFgjb2l2VmryxHQWYDAIhEwANAI2MAXQQ3RK8EgUQSDEd4PaPgItmhJ6F7ywPDgGIEiKp8b4oQYrL65eu1rsA3w/8cTjaII2Q3NIEz2SomyAQmpMBVUpTgxD+jTf9DnMDkFqPO/W9mozQF3aUj8SgGMVAW4BsNSiAfeLpJUVHRDtmYWId8MhWGcKCXihA7O4GfhU0mYCgR4HXSVjBBbVGjNVsE8tLkEpXoLnA/wrCgqaFkAV+RJdDCZ8Tr6vqDdYRpuhEQePZsATVJEo9w30VQrgS0m3z/EOAGj97o0xWtzDxJIBMh3AiFMsx0Ufs8q9g26xtQ1Qhrm7fsiApvDMeO9kyhhXYi0niBd0wyc1+AQYpd9483n5rhml+RoxPtIp6Oa8oB5eHGtNI8MUFTCRpwTAUUbAT14YSgD0sG3Kp3ZmABs107boMUvAPyX8EcDvGKCygPGB/OEugw6g5w5A6w55qsPRcJXqXR9oWFbUtBRBq25vbdt9AeTG+fPna5cvv+L6m8366IZk5ZA5kDnwAXIg7Q4fIAG56cyBzIHMgcyBzIHMgcyBn5MDoUEG2DR64WNPFf/z7/93Z9dWFn97Muw9g+CjQsYAMQ5RRukYwRAgTESq1ZpDCEMoQjMinWZWC+2DFsIXIkv40tnb2Sk2bt/k+QBRcYQmmXkVLKvFAJ8+u6QrQVaq+P2paeYEtlAZVVrYeVangGbDg5VKZYxZ2ujpbnfvl69eee3T25t3Pvb1X/3y+tata52bt7duKMwpoEoSjxgd6VY7gklvGaLMW6bkyMyBd8IBAZo0i9R0abXnVa+ctJutEcukSdIZtCufQFo/DQqwhYx/BfuxeYChp9AQO0XhbQT8K+TbYG1pZumJl2vkO8p9FeBmETNFEbcAMACPKwAG4AICMwn0YKGwctSaYu6DCQhomF9NIwEK04mK+1gNKYGNADQwqRSMMQ+FU52lRlcCQgQ9BLFeu3IVDc9R8fFnnwE8ogxt2YbAGg3yDsAiOGNdxJcAkRpk0plqZ48A+LK+5HNMrSNPraQ2KpLOSIva7JO0pwUtcYI/RAW9Am3mtd7Iw7v3sr9qKplZQCdRl9oA2Ym2zBeB/gsWjUeDAIEEwdQqc9/y5Ead8Q9xkCifvKTTsvZdjbUSHAsTy+i39EisdPMsj6RDMgjsolIcz+YDegoag3ZiJStO0iTekyw1YxQsw+dW1DNiwx3w/YFA1kFvWGyjidvZ7xX7mFsC60Wb9sy6o4+iWtIhPbTreGk+aT/tg/R5Dz5yL/tmRuMdz3s0kY02nDtTDi2wHYuGplv02eTkf8wyAbThiyxpG5I244Fgon9CzOuc4e8JpSuCjDrf34evAmceSsHBLNNbjMdl0jW3VAPzBA23eAcwq+wyl+vz8/P1jbsbI09O7ve77X/33/439a2d7dGVK1ecnYZZy+klf2YOZA58MBzIANkHw/fcauZA5kDmQOZA5kDmwN+fAzMTy2L0v/xPv188/dil8/u7Oy/Wq9WHQqBGGsIzshpkNUzJlCGLVqMdQpSCIuJtCFxqkAlNtdttQLAWZi+NYmFhHkFUk6YBmmUH3IfF0tJ8MU/8wnwbIUmBX6luUCGew9v6aAYMJ80GGStD/NNUG9PpEG2cCcDB+BRtXODQgEeG3c7R55/72PylB89Xv/ud722jqNBFDU6gQdGz/H9MWe4tg5LT2ya+ZYkcmTlwPweS7C0gEb7HWm2WB5owgkCVyjE0pZ7h/gTASBNAQPNKHY8f5f4YQMBRQIhNriu83+au2tAi93XAgGMABJpYtnjXWT8NJfNKgYfDYLTBVNEP7/Eu6MGrS0oggp/wqzVTqjkEyChjngDIZnWZP0AQyvOUgCEAlpdefjnW7vPPfyJA7TFgTYN+BqgV7aIZFksugSQBewhQUZ9t0A8uNcMSmEWkFNIrzSqNk2IBHIE3/KCRZjmDmlih5UXfBaYE2ILuMn12j75aV+q+DIjy8ox9LHgREXyEXzdoC76QrnaY4Jh7l2aKam6FSSV5kvaYYFriqaBfupJJqf2KMEsXeOJwUvaglD8lJtCo7FOZ3ztNBG1JM49+w3dJl57S3FIACHCVtCqAWK/odA4wsdwvdrjiJEuxP8AwTc7LOVLy3XefbadsXz4KVjkuBu/yz7wBYEUsdc7qM16eOa5q13nwQlmX9Vpek0uyhwbZrHjcyvbLOHtonJ2kTVWSvU8x3x9TjyaVROGLbDLeI982deqTbwTP/eZkDGhJlilaZ1UOuZhM+Vsz3dnZqaKRjIrxkelnPv2ZyZ//+Z9P+mj+5ZA5kDnw4eBA+Q/Zh4OaTEXmQOZA5kDmQOZA5kDmwM/mgMK9suXo1z736eLcyRMPDQbdL+EW5qKCIYmjegMRGCloLDpGToUlzaXwI4awhS8eMyL4NFWeQYhsogLWBgRbXFwEEFsARGiFUGa+4aCP9lmDtHZx/MTRYn6xwXutWFyeK06ePjI9cnRxuswzCjkouVIHigAAIABJREFUDozxCY6gz9VqpnZa7Wa93WquotJy6YETxx//xm99tXlqpfXKqy+/fNBBfhvjRocuh7z4s7tODiW7HDIHfi4OJBBHcGBhYaEyGPSnWHxNnPcgyQ8j5L9A2lmE/C2qfY1nzcAuABJdoiSTu3KLJXeVuF3yCB0tMNmPgkqskb4MPIGjfvSlxMgAs9RminfXHaCCGj7q8vjj/BV0EFhKCJGARwLT1BwTjHBtRjrEUA8ADOX4NU3wRS0pzecSUJM0nqybAzSKCcDVD156GbO+neLRhx+hHsETqIQOtdWMkA+ebBiImyS5m/Aa+wT54oVP6UvaSwBs1CGZ8IFian2ZnkA1EoM8i1h3+R7N+a7mnF20LQjQZNR+UVWqz6q4AmSiXwJ/ZIjLeN/tr6BYyoO/rWE/nkdqjskT+UGFgniMbfC9yl6nn7HkzD6JfWk8hOXpG53wEIPANWmnDNFHiSvDjE7GPOqHcrpiZ7igTe0x/YCpzWZZjm9kLIY46h8WBwN8OeKkX19k3Z6AHvnhF068gifODYP8MAR99n8WBPgSsFcpmuzhUuWYmN8fte/iTrvOo3QRQ7oAmd2QpsRv+zwDQem/XbD+mJ+0KXCq1ls5HzXZZDxhlV+46NMOrWK+BYEIviapTJuNBs4r7f5ExLlJG5rQX6PMFeb4PvdV8h1Bw44vdaoDDsWAN/Ci0xl++9t/OX7hhU9W/+qv/qp6cMCZGEGNtxwyBzIHPkgOZIDsg+R+bjtzIHMgcyBzIHMgc+Dvw4GwhUK8GR3gaH9hrn1+abH9xVajdkFhDQGRb/fDsQvyvdIR8moNcxkEoRA8Fb0VpEzgN7QJMKPErwxaZIBa5FOgVNtM7TLAthBElebIUqweWS6WAMSWj6BtVptUGujONFBRqdQm1QblkbHGaI6N0EgbIBwhiU4nPM/Nz7VXKpPRxelwuPbko5f6n/vcZ6/9yZ99q9PrT4bIbIrapWSeJMW34gz05pA58PNzgAlGYD6DLSDqAwI1m80pE3cFhORpfHA9CzChT7yXuV/nrtbYM+Q8R7E+gM5rCP/XuEa8L7B4lrkfA7hQi2wFjR2WnfbGVb2lT9EiCn99gkqCD+SNtZbcLZWT2LjQyAlAJ4FmZpuBGwJFgiABhKQem6eMo1J/A1bQxE+TTGE19dA4ZrPQGfrG7TvFM08/HSCKWV3jAjBUGWUpxgMlAD8ERWYadZFOf0gDXHLRQ1UqBz3qfBJjuQBjIjUBMGpGJbAt0S2wk+gle9AbJYMe6w/YUGIIZf8P+zeL0yG/wIzarIJQAmEBjsELgUi1pSxjsHbpFCALYIk9zPcA+Ui1TXLPaIRWDtSNsvfTFkxN9ZiWxi+qJ3+i3+aCP/BME0v3U/feRCf0ASwNoG0wRFUWE8sdzCv30CAb9EdFH4AIb29kT4Pg2Emv/Y95QlOH/YGWoH92d/+23QRaMj73BctInfUE4BUne6rsmOqzbuku++tYl+Pjnm9wHphPnpb5y7vVSCfvFGPlNBrTESgg7+z+NUDios7YbPF+FRo2iGN4hgLHmCpXWzG++O9bWFjsHT9+bITfy+rOznZjY2MDjbKeMzENYhpGXnPIHMgc+CA4kAGyD4Lruc3MgcyBzIHMgcyBzIFfhANhYilA9vr1m8UPv/c3J778+c9+rlWvXlLjCyEJxbGxMhRCu0KQQk0SphTKkH9CgBL4UiLRR5l5QhDz1DrBsjjtjRP1QobTDxl51AGIaiZFe65Z1JoKoVW0ybBK46eN1hmmN9O5+TYO0BDs0GJrz81Vm81WVd9o+uxpt+eLRqu5jhB1bnFhvv4bX/3K5Zdf+uHe9Tu7NjXH9baaZJS5J0L9ItzLZf/RccD5D2BSWVxaYpoLmjRQGqq2meenQJGfQLvqNFpZmyyOHzIHD7g/xgL6BHmPcd8AC/pbTAdvM88xIZ4eReA/Qvw6kMNJQKJ55yb1A56p4KXD9hHmx3EypmsLXINzKQVA+KFsrMcxYFKAFYxGACwCHFzx42oAiAoQhacEfXCfAVAuBdv0VEHBEOsUVwhAnKJqjrIIi9evXyteefVK8cTDD2NmmbSf3BgEvSyfzO+iAbSzZuALoJ1pXlQYl87cpdVmNMEGQuFK5QRV1EyzXiqBnqT9lPoWuahL6hL4koqRh7zuOwaqBH+HZuoRSOEhaAtNJsCmCeCYZpRqiwmKaVaJFiAaT4kewXt6A6rFvgMoBmTPPe1ZUb995cGrDLUKfeIl9TOlS600RF985or9k9r9oQuSRplEt2NlGcfNh7Hmnox/L04F5vRfTAe7+ITrdDjFsrNfHGByiQJZMbSv0uTlvODuJagX9FCnoQRYja+hDef4J1PZNIekA993xKc61C6Uf4n38rI0r0xms8bbH+uNNulQ1EdbCRy1z44z80oaGWcBwPC3RhE0FukqhwlAC/2E+Cl7e71JXcrUOu7HF9l4HzIbcAR14uomcT1q0iQZYHk6JH+Xkzcrp06davL3qba0tDy9fv0awDLNEchv8DGHzIHMgQ+AAxkg+wCYnpvMHMgcyBzIHMgcyBz4hTgwA8jwjo8gMRz01p5/8rFPnTu1/oQiKpgY8io2TYp5CsMIV+EIHPnD/Io9IAQhJFcRfKsCYoBcOtdGq4Y8VYRpnDYjGHm6nSCbZktqRyi063coBFGFURyJma/ZViDVr82kwp0iFXAHYIgGkch5OiUn9BC0hwjzbao7NR721xv1SveLn/v863/zvb/u3N7cG6rwBpWWUUKKQha8P2Th6X5u5Od3wgHnML7HwIVAbQk4a0dppr7CdYbyD7BSENart7xIXgUYe47nZ5jJHiRxBUDhxwj+WyyO8D1mHq41zP6OczdPgBI8k21cASCLeW/8LASw4HOCVNKd/CwlYAhMI2PCB9BjWtKKkm4BCct4d1lYJkpzF+jQVM+f5JyePCSHCaa5WMu3Nm4XVy6/Wjz1xBOsU5TkSBdYc6Nwf9Bs0XUX4HosPVa5IJWB8gksol3aSMH8guvle1TJewJkZpmi7pSSYqiKOtQao69xCCjv9oX2y+B7RIXvLGqEL0M0rkb4RBwNuQCghrO7ANsUQKgM9iW0othyBHiibsE86xTZs2J46HsVcCwCz5o7pnZJJ/h8SJFpXIKACbiLLOZK4zIbL78Q0MwyxpY4AUq1yATKejjmP8DEsstJwPu8C44J5+HZHmCNcpJVthtjLJn0ffYcYBZ9o0h8cWG8fTUkMCzxgHl3GO+ztab5I3j2Rg01y1qHfEp3AbTZlyT2nz7YXknHFBNfeVAGAVnSuOGzj6nD85DyHdrtQpNscL7vcZrqHe4dQFPVEDFLrswDCDbhgJWhgDYaHj12bHz58iv35lzZSL5nDmQOfCAcyADZB8L23GjmQOZA5kDmQOZA5sAvwIGQVBCqkIIUzIqlZx9/8KFHLp47g0yzhBkSsBXSjOoGylmIYGqAKCw1AMAMCmSeZunpZHjyj6uBxoX1NXhXagvH0AhC+vyZTIZoGijMK9CpoaA5F+ZO3K1HgUzBUhNLBa3QNgOEU+tDDQUAt6n1qlkDbSBpU8G4NTKfxkdZ5dd/9Ss/eeWlH+5fucEhaEXR5lK5IkngluAnh8yBn58DSdOmhWklc7+2sLDERMImrN1qMcfWWUinAcPWAIHG3LeFeABELjL5nkeYP0dmnSO9zBq6TDG1XzS9XOdaIn6ZhXQEAAD/SwIOwj7hOL7GehA0CDdfgANgUAIOrsqZSR+FXZwuXvLF/A5TQeqxDheBOXRI7z0iIl+kEscZs4BYgtaut8jjurN+3gSkKSVR0eb29l5x+dVXi4cvXgwgTIDDk2wFrFzToRVG/YFtUIFgt8FaBM70/xUkzWKjjWhB/2hJa8n2zMcngJ8QkHR7EUUbEbgFvfZbYC/ymwI3otPQgGmg/cV+L0AxATJPqRyhMTbo92I/Ml2trQRsofFEfwSp3GMCUKJRx4RWor20g9AX9iLLmFe8xybLPEGjaeQJiiIfT9JCvsTnxOMAyyIXNPh1RQQ04igzYkwE8hypA8CxPn7I9tAe00H/9k6n6A7hF1sgualTU8uSRY73TONL7TrqjR/qtH39zZmeaE/98MsKwSzngf2Sj9IW9AXvE21T50kkyzOJTbywXoNfgCReypv07N160tRN9aTc0AsGBhhppJqSE/jqRMUEs+a7NqR3SLxLnZrZ98jfkeNYZJ7gfU1HlfxN2sOkX+/806eeerJy9erVitqBQUfZkPc3Nn1/Sn7OHMgceA84kAGy94CpucrMgcyBzIHMgcyBzIH3lAOKDIJHiDcINMg3v/zsE+2LD5xaBRw7RfTCqD9A/qtgA4OSxQTn+SFlIGgp2CD8KoQIZiHfYBo5nwR3SmhaGXVSUEFviqCr2ZBClaCYWhzhc4cIfQJZrY6pwxyHdCMU2jTJ5OmeyRANInD5f1cNoWuEEDpEQGoReRrzsrV2oz74whc+f/W7aJLduLOtJlnIpHYQ2pG5ZpIcFeSQOfBOOBCCNnNaoX1+YaGW/I/VOGm1XkXsX6GOswj5+hg7CmzgmjgAfKgz1x6qV+tPkb4C4HGN+O8zd29yn+du/jPM4SXyLVF+FYCoRT4n/5B4HS/piwlQTPAiUer8TVd6T+sJKkgP0Ia1Euku6TcE34O2w1hBGJaxsbEuBahEPwLQmAFOrscAflynADIAhBy+sVTs7e4W62tH0abjXAzWbptTbsU51OqKCAniSlpjAic11regDdGHQE5sKuR3C+ITEEUtNNe9baa+URsPVhch9o8EVrlvmGaryezUJhNYZh3j0aCYaEap5phAE/uQB4UIlCUtVnll28l3l3UxptH/JoeQRJ2BBkE/459oSjyMdiVwFmJLcneUHgChMvhuiEMQZFQEAS1BI1/sp/F2MIFxbsSpPwk01FG/W6LauwJlnQPMLPe7jF2tGKJdVsNh/Yg0a5CHjr/Bet2jHddDTTiS1GRzrphP8MwRloKSVsvGWFDee0lj/IWQC5Szj6alrZiyEG15++Xd+g3lXU1Beaumnm2FZiLlS35bJurlwUDd+OGr7HPtcPX4QkTQrEtf9siH3X9lmSzzVMXrdGT/0AicotE5XllZnly5ciX1USLKULK/fM/3zIHMgfeUAxkge0/ZmyvPHMgcyBzIHMgcyBx4jzigBISeCMJMUfTPH1vce/qxh5cQMB+dDEfrPYQxPSijyqFMVK3g2St+ELLU2lDmSKAWwpbaIgpHCMN1BSV+RgipapYMMQsCbCuG+tRRwEIwU3iybABlUKHAZZqC7IAT24jhXSHMaO5qqoVAh6aHWmozT+W4rVEqRY6qHqMnZwHs2l/49KevXbn8t1tXr99Vz6yBZQ81hwxJvTlkDvx8HKijUbS0vBzgGCXREqvjv746x4w8DXhyifezxK/opFyBntkPnFa7wKy8JBBF+AHX3zCj93g7wdx/GLPjs8zIVSbvCkL+MpfKTDrR6w+HowYgjtpjrDM+4j4GA+aRKxYehceCJ7wLerhGBFYsY37j1TiLdwq88e7yEdZgcQV9prPiAFzC/xXl9ElGVCzDxbm54slHH8NR/1PFxQvnOFm2Vdy4dTs0rVzH+iLT3FKBqKTDegWq1FQy8BYaaVYaMdGg9Lv4bRx6yR908gwiT2XWYQEp4YKuIJS7dUR/2Yc0LXXfEHifYEYpEDYa4KeL93734PCu+eKY9KCROtRwE25Xuy1MQ9lKoh1oBxMLmuOdJ8dRrTD5Vl5uLrPecEt7mvSb7r0EjFIcoBTxifDIfl8+6zQp9dXdU+DKvtpzQS6nQR9fZD2c9Xv10aplJ6QQYBWX5o+ajdq3ADulzO4QygNSnJ+mC2xFH2gnsshvL/JKq3tx2QdeYw5YF7MpKo04SmpiKviliqP7vvMtykG62oU+ywPNKoMHPAuORdslcTRZBeCi4hr8qUHGkOx7/MHpioVBlYR1ydChDk+7HEB1lzr70Nxgfi1AbxPtNZqfDM6fOz+aazM/b95gBFN/vOeQOZA58P5ywN0xh8yBzIHMgcyBzIHMgcyBjyIHlE78zn+00q7tnD9z4giOlD5Wm04uDrrdonfQQUpBAhrj7wX5SM2MFgCVAJmyr8hZCMnUEMKsHEAIGiO0mj7ANGiMaZNlBcQ8CXOCTtpoqFCGIMjzGARLDZUqLs/0U1NHUBVMq6A6IdhmvQpVCu0GbwheOOwPL0SCFfpRawIUnEL94GS71Zh+9ld+eeOvv/+dnZu3dochKSmAQa7Fo5L8kTnwDjkwN79QWVhYcMqp9YJAX2sCQpwU6CLuIebeKvFqNKI9VkXVsrJK1Q8S70ESt3n+c+4/Yq2InJzh+QFmoUDZGvWsIvi3ucbE9wUSPLUPp+kAZAngMg4QwLmbAjO4XBMRQbo/AT4QQT0BSMRMv1dqljWtpZSHvNQ1mpnk2Y7Lo1wgak49/NBDxac++cni9PGTcZCG617sagSYtb2zE5phHJRRgFQUbX0Q+jMDSqwrLbhETwA/NKgjfzrAukezi7ZZ3ole8pfgjPRFeW7lulfDzMUvIGZ5rwSqwafQGtPpfi9AviFmlAGUsV8NejyP1B4TQFLL7Z45peCNbTm2tuh+xhtPSQNKXgg+mc5Dukdqik90kpc8qD1FSlmf/PRZ3/PeDzkbfE6VpDw+27dZ+eCD5qiCbOyPbr/0dcCeGKdaopGr0361yGqtdoEuXYBv8r40l7VeTUbdm4On0k8Tid4E5qXp6BildkmcgWtpHMgd42K6c9F3J0zZL+mVL+VcFHA0DU0uqoJnYbIqP/mh7uBx8CO1Z14DeUmO/V3TSukech+gWenplgJhrosRfWEqTHvEqVnWRbMMTc1ijr9dbfoGwIaW3cHBBFPL8WtXXpvu7++TnNqIhvJH5kDmwPvGgQyQvW+szg1lDmQOZA5kDmQOZA68yxwIaRCRZXLrzk5x4/XX5h65cOZcq1qcqVeKJTS/asODbnVw0MUAbKSaS/h4CXMZNboQduvK/RClJkETTQIrVJgdauaENB0CFtoO9WobYa0OALZADvz88D5G7ke2RZgdFd0DtT5GRR/NNf3y+w/WGG0yxSkFJ68QYJXT0ChToEMIg4QxfpvQo0j+bI6R8wKnYi58+Uufv/XjH3z3xo1b29SAJlmIiFlikhk5vDMOIIhXFheXQkOq1Z53CjYAsNYQ1i9xesRjAL7HAQa098OReKXDlFzi+UGgmwtiCQBnP+T6NuCA/pSWafUUlawwV1eYieu8rwCSaf8r4lPDHLCN5lODSa2pmeAG1WhqCZAEeFwCSBLiZQivZRQPwMPpPQNaIp1XVkma+feBE5ajtvRpkagPUMY7PwCCxec+/ZniicceL5qALNiTkgl6PD6RGnUgPwBwuruxVeyzXgVjluYByri7H4h6uf6TNpN0AvbMgCfT7E9q036oVQToJgukkdyWs6+pD5SnjLtMqbkqIEYieTDNRnvMfcLTKUeA8foslLYBzwcH+wBL+PACOEtQjRpjAlb4LwTcaQgg2T51yzeGO2j1ZosG+eooCPrcH0J5lSz2yx6SkQtu24eoJ+VGn5B0+2/fqMua5ZH5AmBiZ7KpqISPGC4pkk9+YeChCJWiD9A36HOaJaaWPe61ucWi2p6DNkwpySsA1ffLCNvmCrocM+qQn2N4Fibv8FLe2bZlBFZtOnhtm7wbnEbGJ59l9JEywaMZGxyuCDZHf+yC/faHOX9YTn7bjmMuaGY1vstO+hhcZQz4QYeMsy/gdwvAsU9VG7zvkGCLqGdOAaGr+4CA2P5X/MOguaVf39Qpy+KcLOifkiMxexsbd4dbW5s2EGQlQvNn5kDmwPvFgQyQvV+czu1kDmQOZA5kDmQOZA682xxQ+FBcG/twsL3fefLi6e76ykK7Mp6eBnla6h3sV/q97qiPRll3/6CqOVMPYU3tLqUdhWaFQrUoIgCKKWSpneFJloqGrcYSQlqLvPNFt1tFsO7zTNqoXszPr+AvCAL6+CdT0EXIa+NbZ4hgq3ij0GU7akNIqUIbUi6CZiRWORjA8+xUDRkgeDUQltYQmx6Yazcmn/rUC1vf/OYfb+4dDAYIUsp0EknBVA33HDIH3pYD9Xqzgt+x6exk1iYC+DLz8TSHTzzE6a1n0Sbj9MnpLnF7aM40maYPIKhfADQDBa7cZl38kDn5miAY4RTPp7irYXYEIGEd0KFtGnendVPfY4BAzs9YQ+Rl3ei7PJbADIDwWWiBSC4BnpQuiOMkjxUSeWLNkBjAmuuVIDhh+UMgJJaDKcRxHTt2rPjqV361OLp6BO0rzaPxl+6ahg7oi3I2oUYo5qBh+re3uxObyLG1VYBtQaJUW7QLTd6t3dWrT7D7g+BNdJ/63EciL/TNABTS6B/vLnKXuXQIkHl3v1CjTHNuzUON29/vACYdFAfcw+cYeYWwqDr6Dl5T1KlcEMd23bcEi2Sme5YZ5aOAWNw1xZyl3093gEJWWuYLIMxaUvlUxuSkWUXOFOSN/aNs9DvGz1TG9L7n0MKirKBW8IgxEJjsdjEjpY3hFMyoiSsuADRcMWJOyuEDszER1EMDK0AxG42xpk1D2S/pc35Ih/nLYFvR79k8gahIClp50tQ95UnzKZVPPIxy8MO8jaYHtqT25LUgqiEBlPadOUE+SgricZxlDe1MGsVkkvXFmphoWtmzBpJVT6xTP12Z9Hj3xMvQODOC+HnqP2o+TrXco18HV6++Hs35QUidSM/5M3Mgc+A95kAGyN5jBufqMwcyBzIHMgcyBzIH3poDSSC5J9y8da6fGetX9IovE6T94aeeeeTG8ZXF1Xqt8RzaGOvYeiEk9waaLe3v7tQAydD4wpxJgQzhTZkmPBDp7AuTKeTgEDQVhDSjrExxJD1Uvjla3L7eL66+ulds3BoW165sFTubaoyBDNTmiiY+bXqdbpgS2ZZymYKtspsmm2pJICvFaZlIaTz7L1g68Q1hUEfOceof/miQAasryE3ncSRe+/Wvf/XVb33rT+7c3etiqqQmQvwkVOHvYI28zeEfLQfANRqVtbU1lLkmgC771WazpZ3l8VarpZnkKSAOhfJhvVLv1iq1FoDVaeIvoEG1CCqiGdgrCP2vMYsQ8j2pcnKWKYXfstoxDrJYQzNnFbCoJahBqPBcEXgo/TSN9Kcl8CO45GJAiylpXiWgB1BhNjgCMoIPAheAUCwYViKvxNGgz/4IgtgX8xlUBktNJ8BGH1knT54ofvNrX8OMGsfnAOKubxeiWlgkR3nBMkE486uxJDC139ktbl27ViwvLRZHj6wCTLk32Eqi0bL2DYCR6jSvBOAigxqoUpPi7mmNufZKegVQNI0UBAuTSnmEeWYc/EH9gPdoi/WLvb3dYmdnC01UTnsU1INu61WrrQbv6ty9eIwgTe5d8k6wUQBHPjE+iWrZx1W+m09fi4JoqZxbieUtnPgvwBfvthANkeZQRIvy3hbSm62lp9l4unFSJgBO7+Z2jL0sSu4BpugD+n8w5PxfsNn5pTUuQEm+UDhAA3cHHgzYUO23oJ88to04YTT2TN6i0XQ4ge1pEpnmhdSR366YyaZnEySlO4dIJD4BibP+8G6ItNm4lWCYpxhbvwCZhwaYR61i7x7m4lasDzsDo1wRHLYt+u03K3O0gxvLyojyVcotEgcBlX2uAQ+c/FrB1H6ibzK+r6mtcjXgXAcNyL2XX35JyuztjEKecsgcyBx4XziQAbL3hc25kcyBzIHMgcyBzIHMgTdz4FAYe3PCz34PMYlsyoZ8PV9MEFOWPv7IA0e++MmPX5yrVZ7HZ88nMKVcG3vy27A/2d/drezubtfUKtnZ3g7heILA1kbA0TRSh/xIVCHPKRAp6CDLIXguIFAtFbtYvOx3akV/v1F0OwpUC8X+3rDo7Ha5cyAAQt9cax5tMgQvqOp2OqFt0kYTAf0V8LBqoWtqZR6fAbviLhCHFg0iFyIh/si4ehRvonewQvyR+fb87fnlpSv//o//4iDkTGpXGouK/g4+ydtfgL9/R8056cPOAey0Km2c04PLVHrM94WFxSbvK8yHM8xtgK7qkUaz6XQ6QIgXUljjdhrBHvCLmVgUN3h/mfhbCPFgtlX9kZ3gvsassh4A3PEia6QdQBHrRu0sQCS1ZQJIcpq6hrwMAZb4wLxUa6ycm55mGFALcQa9lbmoBTHKsrRLCrkoaz3e1UYy+GwNJ06cKL7y5S+DIKOKidmkGkmVAMMCsGCN68OLMlwBdrG4BdDU4NrbBpjq7AGQzRXH14+EnzFBMOvmN/Jb9n56fDYuxae7gJnAn0CgbaitKtij033pH3IHqQ/+6LS+D5CuGeXe3k7c74Fwgm+CQ2gyofFk/92TDNLke+KJ74wXYwa+nuLoIsAmu0la/6aHlhlxdka+Bn/9AsA8jnf0Ux6n+uNuGj8CfdbhOBti45Ep941h8JUoSvNjJsc4Hg75M9L3Gqn7OOnv9AAuGwv8rhRrxx+gb5ivU+bOxh3m0QAabTO1q1njDPWK/hkfPIbX5gNUsiG00KLleFZLbASCKl2pnqQ1Js8O32f9kSaDPJF60w0lv+WXcfIheE6/yjzyPPpOFHcvzZIde271JfLNERWM5S6h7OuVOaunOlUr+3aCgHnyKPxRcvCLWp+0UQzu3r1rHoNEJcLiNX9kDmQOvJccSLvte9lCrjtzIHMgcyBzIHMgcyBz4G04gODwNilvE62YEN/Eh8QwVurgqn/puUce/Zf/9Dc+Ux90P4kg+rFxb3BKU6ZRb1/hvTFBa2OCr7DdXgdNigaaX/uAWoNivtksWnPz+CkaI2QBtaEZoE8ga68UraIxj5kQso3yVKO+WLTnW2h4NJKZZquB6dQQwXcMUDYt9nb2MMecFM02BOJnDP2U4nr3VnHkOFZpCIjt5UVMizD1osvVVguBC40PtRP4QctNwQudiDFqgoV3AAAgAElEQVSe1PWH1tYc6IH+/sGv00qHf9j+L0i4pZgJyxS65ISvbxmoKIS+SEw8e8t8OfKjyYFSWv7p1ZPk8YP9fSZIrXLkyJHG3MLCHCDHEsL4Wq3RPObsY90B81ZG2IatIPjPo/4yBAzY9Vw+ELEOEM028SyS8SLTso2z9TqmfWPkeZ2Oa/Ib0FYJGoUDfEEh1zPz14MrTJPOAJNmbA7AKMCVRLmnulrGkw4FdQy++5NCeU/ghUCNYJwIgg7kBceW0UL6/Gc/FwdlaOI84XAN/QiqubW/3w1gQ4xNOtRGIjHAKwGP7c2d4u6tm8WxpZbrL+pW8600uW420RQiXpqiPKcWCmSVQQ266DMRofkUdKX8wEq0bbuaVdpm4o/l9TE2QFMt+s7eZBtlvQFqAb60GpoQws4YyQSK1RqcvkilsqoEkqSlpAE8h2cPGWHXMB+bo7uK2lZyN4CgkkYLEiuYJRhnfuuRFjP6nN6JE6gyNzhmpM/qiEg+BCzV4KKIlQVgZ9p0CgZEvXOcHjpoT4olDkVYXhwAGraL1uqx4uLDTxQHfb5cWDxaXL1+K0xMx9JvJdA8ZN+0vUQTG70djHoZK0CwRp39lj1cXjbg15AvKCIveaJc9K0SfvgsZ1yaB+lLEMdP7TBZZF8F8jjZNbT40EgOsLGBdrBBM9kme77jZB2pLguSyOW7c1OQTG1D+n2UuDp5/TMl2IVlc/Ukk/0Y7f4pRbZYc4DME00ur1J2DtDtxP5ep37u3Ln+nTt3BltbW9YLeTbCR9x8zCFzIHPgveKACzaHzIHMgcyBzIHMgcyBzIGPEgcQRYpKAxkOzbHGZ559+Kl/+y//+dda0/Hv4ujlq+hSrE9GIxyS9/DtPESRY6RUpdyJNVF9dmKdZkv4uUGQQYTlF6EMqVMNGv2SVeLgPYShocLiHD7FEOTVU6s0Q+NhACjWbOBkGu9nY4QyzgDA59GI8s0ZOABwNk6mUgrxdU7JUxNCQVMArAFApoCvzJOUeEIIJUMVP04Yd2L+Vq3U53g/tXZ0vbvf3fvOD//21TvKR1xqIRjuSerp/fBTeM/fCOX9MDU/fNQ58HZDGpPcmVapVxaXl6rrx49jPllZQ6tI32Pn0C7T15HT6ABhHB/29TXkb9yOVe/wvkW8wvo++MgG9z5TdQkBfh3QbIm0FvOKiVwsoumyClAwN8aUchQmg87ygJ4CaBAsEkQ4DKxYmwV/m0XxPENTaP8NeX23shRST8s8UWZWh2aSzfZ88cIvfbI4cfwE63aIhucBaxKTRoAK/YWNuauNJbJg2SprTi0uAaptNElfv/Ia2mb7xfqR5eLB82eK40dXI6/7gWCcYIhgh3dpEEDxWSDEeN9Tus/Jz5kaY55C2e9rPtkrel3MutEYs03vPdrrQ4P8ETyL/s56q1mfoJwqRgItarZ6ZyzSpSYYgfFIWmO8B1DGvlLWo2aT/XRfMc53dpeZtliqR/fyKZ5BI49X8GfG27KuMo0MafwcZJ55iXef1Zgz3f2VT6gzL/PB8WUimUf+C0axTRYDDhXe6QKWrZ4sLjz4SLGwdIQduFagMVVcv/oa/UxtWFMclAIvPOTBOulR1OeIeoJp8AEUMJm0OkbmONTsSsBkzLNEr7wLeiIuPRvnWBsfPCGt1Bgzroyvq3VH3nIsSn6V85x7yh2IpE1PIK+qFpn3MXW31QqmPkEzAOpin3hNLA94H5BvnndAtWqD9bq3tnZk78aNG86TxED4EARQIIfMgcyB944DGSB773iba84cyBzIHMgcyBzIHHg7DiQ56u1SI74UTu7LFNK1YgL/wGhaufDiLz3zzH//X/9Xv1EfDX8LXY9PtNvEIuBwEqSCTBVznEodOyUFn8XFRTS2FBArPC8UC/NeONRHiJ0AZiFN478I8xakoFoV08gRgtlILY42wu60OOjicwwQTLNIpUG1ZLQJa2Na2cNJP3IPmmgKuDj0r5CvQVuY/iA642sHfAFFBMExpFfSEVmlhTIh+GEWRAWhsQC6MaTvqsng/KzaQsus84nnPv4XP/jedy5fv70tnAc26MEE6snIEt7eJDkpyOXw0eGAI+j1TsO9vE4o35hPzJ+Q+0FXl5ZX6keOHkWmb6CVUj+JL6UH0Q07DSbT4LmPe6QJ6iyY8U5XAFJ8v8rC2GBGinYIR3RZPrjAqhzjvsZcw6dSpY0Qv8x1dDgYrGCajCaaIEYCHwCOXDoK9GgUJS0b1MyCpqALOs0ghOH6SWCGWku88hGFnc+8RznyCeyEOWWgL4DXlmf9qXHG4ioee+yJ4vEnn4RqHMADjo3QHlNbVOBbcz3p0B9aAkAAZnb19bVb3Lx5q7h9+1bROzhAu6leXDp3unjs4YvFkRUU7WBpI1AafV0lDbLAsqEmfFBxjx8AG6AZegzLBAQ12fSi/2pxhd6Pz3RmOMLUmzTzwT/KyyfBMU7IRYvO0zYF7JvNBHgFOMa73Qa9lHMB3lhQUEhNMMYlrhqHiYRJJXWWWmXyNp7pi3sf4xt55J0wk3fz8MFvuqzv/nD/u2aN5osc9mE2HmEKCi36mnMAPZYx6qR+jA5nfYVoynJoBCBdo9g9GBZbB5Vidf2B4uFHHy+Orp+kW9Via2un+NGPfkBW+SNNqQ+OpVq/Y0zhQxPPsSe/6foZ06G+Jwc7caJPlJX2GAd6a22J3wmwNb4MkHUYUn8TLxwn+UeFCTSjjICjYxfrjCqcG+7dhrI9Ske7Oh9jnGJBMq51+LNAlI7L+rSvQ3/fIaxyB5q3Gb8F4tHuDDPMLgV7y0srw6Nrx8bXb9ygEXpgJ2IEJDpejMghcyBz4F3mQAbI3mWG5uoyBzIHMgcyBzIHMgfeAQfuE0zeQe4yizASIlaBDkJRfOKJSyf+h3/3b78+7e7/DlLw81oBIWQgmU77CkwIITU0tSqtdgtLMnTLEHBwfF/M4eMFZ+VFCzBNh8yAAJTDHAu/YUO0PjhZEn9icwimOGiutdHiaAKQ4TAGEAyJCQFJOQefYuEpXEHMdhWNFDoFz0Ah0LVpYKND1qIxB2hXBTSgHQXZKhohFQU6OqOmh4JloyEtCFzWXKuj9TauIZRGJoSyMb7S7n782Wdv/cH/8X9uqsACIYiGFax+ELNCYyELTOUk+Sjef97lEPlDui9LJmmeGV+snzhZPXrseIv5NAdescy8P42wfh6+HGGyGcB4a6vc9SeGIlZlHxClzx25G6dJCTADpMXReFE9gpw/R4og8wLJJ9GUOo1D/UWea2pTsebCQT/vILbJx5cYhmvKSR718kR6PHvnQQwi4hwveyG4YXlBljKvaSm44gUrMI1zqtPPxaWV4pFHHi/mALrpBdc0tLO8q+GlFhe0BTA1BkDbxc/Yndu3i62d7QDKejjyr1fGxUn8jn3iuaeLB04fB6jC35edZU0KetgmWE+AI9JRmvhpGm26WbySY3ed5EMjaxzVVbMHTRPMqsu80qlyqmUEwQTH4plG9KOV4tTuKuunfTIIislH09k0olyZJ0ChoCNphemDTABMp/xBA/uSZRhB8Bj3qFRnpFFvjEfkJAtp5XiVd5NkucFxSuNHgwaBJMGwtHMd1mUefs0Q9TkOaC/GISYbm51ip18tVtZPFw9eeqSoslFO2NE7jM/lV17mi4iD2CdBcqNd/ZD5RYKNl2aq+iyLPgYv9dGmL0ezpP7FXKJN2y2DNCWwcEa71AWdqXdpvB2be/z2WT6o2WeINAFH5qrxQRt51B40eDIqdZLi0OOtv1aXLL/QWGRuW0QT5QYPa97p4C7FBsSroSkAzdkRA9ZiUYP26urq6oh5OtzmAAfaDhzZduRrDpkDmQPvDQfSzvne1J1rzRzIHMgcyBzIHMgcyBx4RxxAgAjh620zm0H5lAvcafTip54r/tf/8ffPVof9f1adjl8EEFP4QCYf4SGZI/yQWBFeKpoy4lusMr+wVLTwVYMsE8Ksgk0CpZLZTAsBCFcwRRfhbPPurdBAaQGSLS+uIARx4hrlPf3y1o2NEI6Q4ND2AETDpHI6xlsZVHlinAKUp+A1F2inxVFmCwq0AAUAZGo66JusqCF8KxgjaIX/G4kiqEXREP5T9lHlQxFMQaxabaMRt7p+Yn3wlRe/cPnPvvXNzm4H0zYEL0sG1EDnDTIhh38MHEgjX/YUYKx25Njxytlz54v5+UUmXbEIDLYKsLAGkHKChbFO3DygbwOQAI2w2klO4mN6VdFgKbpMuaNAWmv1al0Tyz30biaUm+d9jvcJ03CEFswyOlQXR+PxGbR6GoACnHMBIMC007m44JZAAUJ+mCFqUsdjgBRqfAGVxI8z1ksw2Tz6tUI/JwFfkSb4UPYv5RUgEUweCXgAtMwvrxTLR44Wx088UKwfO1WgLYeJ3gYAN2sY/4KjMKMEJAOwEHDZ2ekUdzY3ANA0exywzruss2Fx5viR4pknLhVPXLpYzLfrxRw+vqAkgCi1wLB1i3XquhaOBhqBNqgHqnftqtAj8C6A5TIOwESQTQDNPJSP/HyoUOQBBZYTqBHAEsgPs0rBeHxoGS/wJaZlG4JaAOaxV9UB0W3L+oIeyrqHBOgugCRt1hs0C+gI1iWgTf4KULm12IZjEe/Q456htlTSmHI0o6YYR9NiTyHOwPhHejxbFkIDCJUo3jQytA2RnMjD+MYYA2hJ+BCt2+1Ov7i7PylOnn2wOHvxIcxkF4JftnPltWvFxgZ7LLyqsE/yAM9sFfqg2+F3fkXdjI97pjOrgdausFQAcZQpfdpZVoKiHxRKJVMdkqQGmrwkR9QZ4+mbcbN2vFuPcf4NsQ0FaEswGvQ11Wu8Gobe1agzP8+hvUz7UzTJKvhUQ0W5wCdgpSlAxp8rT5edp7UJc2WXQeCUS6ocTThrplYdjUe9M2fO9NWc296+q0Y0yWUveMwhcyBz4F3ngOs7h8yBzIHMgcyBzIHMgcyBD5QDM/HkkAYFmjcENSBU0EAmQfQb/Ze/97vF4xfPPj4d9P5JtTI5p/kSgsZBo1mvIyjVES4xrUQrS58+LcwoEZQVLuoIwAqpmkki6COrKNii8YFgXwHEqpK2hybZxsbtorPXCW2z+blFQId5tB+GxaA7QMjuIQApP9Uw0cLHEdopOvVWm6YOADaZHiD0TXDoj48kQLJKjfgmopRYWZh4IkDPhF2FRsUdzaQUqsdqpRGJ0CcDVMEZI1i1ELbOaM5z5vSJq5ubOz/5/77zQ89Ho3SVXiWRUUGvFB4pFyEEwzfzskzM948sBxKApIxeraFBVTv9wNnpysoKU6laYw4sIVsDeBXHAYH1OcYpEdNlgJFlzSq5HwVs0o/dXdbEFQAV/CPhPLxSXcScb5dKMa/kmMFp5QgYM7J7BV9krLLJ+ARlHsS315FBXyAM+R+QQhBAEERgwPnn3cDjvTCbg07qmOKQbj4vgRkN4QTMLFOufevyGY98rCHWF23UGu1icXkZTdAlkPJ2ceHCo8WTT3+seOrpZ4orV14vNjkJcXdvL0CxPqbTaot1ML3c2LzLwRpd4ve56/5pXKxiZv38048WD5xcL44sz4f2GDalsR+Ij9h2MqcWJIIwftUqbapNBFjmvqEGmMGNyfVbrjfvgmXeARm5u8YTcBbg2QwYs37XbYBpgl1k9HI/ML9gVwLbEpBv24Lr0iFwFppz5vE58kM4dAlUCSj5TEK0wfgGkGe+IMjdj/Rokz6ktkmbjZt0lUEQKoXynsqxJQWNokSx/5Apxo2xK8evrF8wandvv9jk5N8ObiFPnbtUnLlwkZGwHS7GeQOQ88rV19gHUdmlTvBc7vKRLyQY7+ALe6f7tft4AqSkyfaTmar7vHNGoBFNR+aW+33aGwUH5ae7q3OPXkS3rN/91Xf5IyAlwCXt9qt8doJGf2gy4mOs1F5LfIn2KGvfuZi86OylcQUzwydZrbZIC3zHM/UbHcwqpychwNNhp+Tbwf3kAfF83VNdBGxmlk0FzHqXLj1U297eaezs7ri4ykEI2vNH5kDmwLvLAb9uyCFzIHMgcyBzIHMgcyBz4APlwJv/41fAeENAuCIcCgdLSwsVTqk8waliCyNUUHDKH9nr1SZOx4YIRwBgnEan+KMPoNYCZljtOXyI7RdthE99DzUQXPtoklQor7+wOr7GDEvLc8V0a7e4df0nmGTdLB566Onikcd+CYF6rZicXCiu3+jgZBsgDbOX0RDBdaRwWsds0zb74WR7POyEzxxNvRoYqgHBBR0Kdg38DOn3bI5TMaUTx2T0jP55KdzO+o6gNBXYMyQRcvrk/u7+r507e1YJ/y8guwM0oUgXgBoCWEImLJDkvhDUfM3hw84BR9hwbwjTe/qMecxjMuENubs4dfZM7YEzZxs4N59ubm72nGsriytzgCOenrfO5X0JQKAJTCPYiu/3Oo7J6kusr03ebwMqbPOsRsseYAmmXdMBvvGAdouTgAZLAAOaX056vYMltLdWR4N+K8wqnaOAA1pRqhUUYApxOk7X/M1kIAuAI2Z+xAkUhxoazapZQ7p5yDvkQdNF+zjiOQEXM7AM5ElQe8TaaKLR2cIpPz7M0RACMGnMF4888WTxwqc/W6yiUXbltavFH/7B/1709raKCetP73/g5bEGBIJcV/JITq+vLhVPP3apOI555Qqny9ZYQcHjWfuiz/Zptr54xs8XfTGE3tIMPFHTQB9hU7WzKJu0svB7JnIkOAM4TtUF8HcA6GwCUYf9TwBLApKoLt7TSmc/Yl+wPoEwg34N3Rv4jbv5BG30W+Y4eAV93APThNeJXisu0yGEEPwFTHLXAJaJOAG/SKXNCDN+lftICcnAlUgGyIn6pbv0wxV8obhAmGak+lusykfRKOqXc9Ld63li7xxO+peoPmmFqUU3v7RYPHDuXLF+8kTx2uWtALgExPj+IXyzzc3NFatLR0P7b2d7o9jb28Hn3AHtj3jejzk1RsNLX2fNpl+K8OUF/YTxoVEmGc5P4K/4QgMEMfhsPoie8QsS1UyD7lIbUsrlmUCudseGGprJ9lHuyWdGi/HAftLB5jK/PtMEcfucUFxvYvHMWGFbaXHUlaeYOxfL0Hp8OOwfgZClCcrPMOQvybcLrZhbTqb9fr/OeqtuboOsLa9AAjM1xuit9wkrzyFzIHPgF+PAbFf8xSrJpTMHMgcyBzIHMgcyBzIH3kMOJKkE0YWHsf+8/Ke/9Wun1pcXfgnx+1PV6nRdwQ3BgsMnlbQR20LXjEeEkhTFHWFZLQOvFo71sUpDmCGrWl9BPEIODTTxTabT7MGgW+xw0t2169eKg85+aIKofYCZTLGLo+87dzZC6J3nQIDxSKANMKsyQKDvI8gDhNUB6GopTmf9CmGaUSmKJu0GhSrpTsJ1EohLQTs0Hux3/K+mkMbLPPnXz52/MLp64+orL73y+oYZqAXpWTkNtCw9eMvhI8UBR9LgSP90MHUGjoX12jPPPVdZW1urdbu9SrfbnzQa9SmgwEKtUQ9gDEAHn0aVVdbEES4wk2oXv1lzWB+fpaol4u4C0LzOXAQYQ68FJIb5gxlYAwKmgmpHicdQuPDEvWW0x86iHXNhPBoeQ+slnPMjuFcAEYI0566gUFKakf40M+2NYIoLV9BAMNi8Scg3XwqCadhw8hLVpUgAB4EhzaTnFhZZs3O8zwGAGLdQrBw5Vnzmc18slpZWA5R7+NFHihs3bxd/+ef/QRwGc8sBQPYgtUfbAjk1wI+Vpfni8Uvni2Or88UaoMzifDNMK9k+iiZAVxNTaLW3YErQIZAlXQIh5eU4GS/IFM8zQEr/Y+ZReyv8lNEdn4mJOjWvdA+xDfcagSHf3YvcC/R/6H5l+03AHveGunmpV3oEzNJ+RhnSyv2s1FYLWme0CNYJjhmX+sBmQpztlP3hJeouQa4E8Jmcxqgsd9hvZ4fjRxYDvY02BMdiTEkzb4ykfHD7Is4Cah2qQXb15t1ib1gtHn7q2TjB0j3aPdWqtra30N69VWxu32G7RKsXYNFaoiZAr8cffZLxXuEk0gQ06mdOrVvpGcSXCfgLI1/wiX6q3SsoBmQV2mb2RzqTSey9uRhjRtqhvzi07pyv8jzS7NPs3fKOmfF++WIeAVhDaPURL4hsemi6hYNKRo1MXHyXM+IJx5bTKjb/lSYpaJKNV6m3ZTNWQxNY91b949HhsIn9zn7HDk886RM6EkNtMIfMgcyBd50Daed/16vNFWYOZA5kDmQOZA5kDmQOvGscSNLHrDrEvtrv/favnz4y33we9a2PVybjNU9Hq1SR5fleH40TFBcQzdS+QCBXu4u00ESp4xC6hsAZggzCqlopzXYLsyUEToVXBFYd6C8uLRRzmGD18FfU2ccsCMHk8uVXijs3bhY/+N7fYM51GQ0FTs1DE2w8xtl3bYJGC37GapoGYWLZBChrjtGW2KYtyFDTK/7rEhxDMEPkU8BViBI0C5NLBSp6YByfCn1K295HCGFIVaixTIs1hNfKl7/4ucuXX/7hK69cuSVCoZKGUqJyYg4fSQ6UU7wcwgRiBGrANIipoJ4KovVTzzxTW15ernQ6HT2fDxGkKwuLS0vM35MAHCeZ24to3tSY+hj4FnMANSPM8vaY43OYpJ1mTi0AuGwxXe6gTTZAbG8xp+aZX3OktTEbbCO0A7p6auVkFan+LCdWXsSM+VR/MFzA1DHpAzGJEdU58hKwaAbWqEujKaQyvEAC6zEm5Xjku1gJfeESkLFwvJIgACKYo7aZgJLrcG5uvlhdO1a0MXEGuCOvPAGwwCdgExPLpz72XPEYgIkmh1QVAMjXvv71ogsw9u3/8B9jnY3xK4hJaPj/awGELy/MFafQGju2ulwsLbTj3gQYa6HV6eEdTerS3LHFfiDBag25gNlOaBcqBZSIw3tbxBkfYJpAlHGsbcGScCHonfzGBYhC+chL3a55zMFnQA3xVKSZpGW9apgRBk/hhWVTeemALuoUoGG8RLzIJ7jG3LB94qPN2HSkxU2HeCaD5aSdj4iT38nVYXqNeAYk6i2zxdyTFbN5Obv7Zl3W5IcAZ/IBxpjaXmx21g+dPOsTrtfrF7u7neLVqzeLaWuleOyZj6NduxBO+gWUNJc8QLMXMKh45ZWXgjbBVXkBUbFHPnD2QvHA+YvF9u5ezJ0mGoUeTMEH+mnMNibCEC1dwVZplG+aPQZ/eJc2KTT4qbZb8MSU6A98Io/P8iGlkc85SpwgmXd90zk/POzFd3nufu78QROMcbBdNNec47YDX8lm4M9RtYJvMaHVgIuhiMGbtklukd9TZ/mDxIqcTnvEHbDu9u9ubh7s7m6Pjh07Wtnd3dGM2rriw4ccMgcyB949DsS/au9edbmmzIHMgcyBzIHMgcyBzIF3nQNJaknV6spr6Rtf/fz51fnmx/FM9DGEhWXRJ7QzxJVC2gxhJoS9JDyqpdBAIwNZCUGMr+fR+qoihCs3KlQqjKqpkQQxHD5TTYvT8cAdEPCqnHq3U+yi3bC1tRl+jjTr0VRy0N9DsFa+6QGY7aIBAkCG25hma4RAuINQNKLNfhKObAuJRzMytWF8UYBT0FKAUyDTL5rCr+ZgpmnmQ1CrwIBgpGA6mcdJzfBXfuVXdv/k//3m7e3dbo+iiJK6////2XvPYMuy675v33zffTl0DtM90zOYnANmgCGAAQlIBBEoyqBFypar9M2hpCrbH6wPLvuTZbtc9gdXqVQlu6iiRKtcKtsq2qIoiaZBEIHAEIMwAKYnp87p5Xfz9e+39j093SBAECI1wABnd9937jlnnx3WXnu/t/7nv9YWaSgNp5DWe+pHtp7fGTpt3+KaHXFYUzpw6HDl4KFDld3dHdElcSHwq7o7Uh7lc6xea+FWSXD+Rn0WoMsNK64wP3YAShbMwwO6TXZxd7yGDb7N9wkAmi6XS7CZ2uggJEyJmJUOQerXOD+KoX98PBodAGggLtIIr8kcD4xnQ3dtV+gxRxskiCA4IAgmOGFgfXsTIAoKLChBq0Op3VVRgKvO3GzhAt2BKQbYh5szccaI++d15dAHdMB3GpBkhi1s62n/wWPpbuKOre1z7wHnEcxLjrp3fuQjz8Aymkuf/9znolZFJyTNNE1zAGSLs600126kZUDw2RZAHPOeTTAAySifcmDjhbRpInMNwIlSBLnC9ZnyTcEUE2DiVBaZQJTfBbcEawTTAjSZzmufbwp6IbMAyTg3ZVBsCqBxz/vBHAugK4M0ylZZC47JIizqCnAMIMZ7Lns+65oSeQESPZd5xlhyORoaboG6uprfe8rO5O04RjnvaKF9mIIx1+/nL4KcStxyzS/wxNGxjUQd8aw3ZW+5AUo3Xb26nl545Y20wOYK9z3yflwQDXVnXk3SSdoGIFvfvMYLiUtstiArN8vG8ukccR2XkhtROM5uuABCHGu5O142Aat0OVXnZJXtES8yWkPnvK5cjPkWIBd3PIZcrFm4SiFwyGNEfs792E+veSy+m911Ouu5uxDL7Mt5vR6uxpSvcKxH4M52MfZMWqeX48Vbk2gg2ewc5GVO3c1ylpoa1OWLkT5ldDuznf7sbGcIIFfRJZRNJnzynac5KVMpgVICfzESKAGyvxg5lqWUEiglUEqglEApgVICP4IEpiban/Uv/MIY0EoSIGt/+pmn9q3Nz9zJLnD3YEgsupseJge77cFXICK+7LEI0I+BrXEaxg9GjmwDDdABBpvAGLSxbFBiaMo6a8Na0aXLXfIEzNqAZGsHDrJT3loYRJu4XLrbZQ/3y+7eJoYXwaLHxBsb+h1bBnBsMsFwG8Mqq08i5tmIumyChrGMAtsWbA/bg2HobppCHfbB7xriYQ5iRGkIanRzD/ALQysbVx2M3P2ddmv42c/+8ktf/sIfXL54dQvgLekf56MFoPYjjEiZ9ccrgULFb2xFcS3UPlCZe+67t2JMI3QIws2ImPKtZQCTY1jat8AkWslKCXEAACAASURBVEO/CbFXFwzzs4kqvQbIgOrVHwSMuR2DW5fK15gTV1EtVL7W8jn0aQ3WSx0G4y5HNG58kHl1G6050usRlL8/mIHJwvQCKArD36Pt050M12HAG0EqAV4N+CEAcoAEgThobkz7YD6YWolg+02AsMWVfWlpdV86cuxYWlldSQvMO4FsAWMBDd3y2Cwzyu7gWgc/lN0r19LawUPEYDueFuYXALfazBHmL/+sfwdg5ec+9JH02V/7tfTcc19PF86fw89zkDqtegBjHUCxuQ7108t5ALO28xwWaVN2Kc10fTAAvL1zftpnwSTBFfsouGFsNbvkobhGdua1QL0sL4GWDEK5/uhu6Zw3r3G1mPkckQsAkOA8B47UNV2r7E/s3MlzfhcoEiALsIxyBBW5EPey22TOw52cd1oO4x/tVTa5H3ks/G7jLdf+5KOrMmsP57EGcSxSzkM+O2ay3Ol3y1YVIrB9lBWd56qujHzHrbXX2yNOGHEdL15Mp195M73voSfSnQ8+Sh/wNERmTUhTgLC4tffSDhspXLh4IW1tbkYblZ0AmmBYjTE6fvxkOnLkaIBbqqKs2x47BzteLVxwffnQ3UMH0cten3hwgKtu4mI7BMpwZ7zeNgFK+xax3BQWcrEcgbMCDLO76qLXZTL6xW45D8zjmAiUCZIpFcc4xpzr1m2eYhys2xcuuPAz/VJlgJsysvZ2CJ6yDIQ5i67NkM+NMQh7Vhnwe27Sbs1MGOvhoD8cXFtn+t4wPjxTplICpQT+giTgKlmmUgKlBEoJlBIoJVBKoJTAuyoBjYRIf7Y/8rFHIyOEr8oEM6T7zKP39A+vLR3HrngY639VFyXMFfZGq1YwmGsYHhhnWp2aIRqAGkIao/7pg7EoS8RbGJ1+8brxjqoYx3iYcQ1D13hHAFZtDHB3ztu3b39aWJxNWzubYfBpD1Wr7uK3l2Zagl97WE1djMUcj0wXTOPoCIzViEEWRjd1GrxaRptGlLvgFTumaYx770bjNNzVtLowI2GTySggojSBeaqVBR6sd1qtt2bn5179V//6S30sLoOQacf5KdNPjQSyDt91733EBm/JIqxinBMzjN0oq7UTmNfHUcQVvhMJHFimUh0BgLj73Rb3wIFqd6M3jzCFOlx7ieNLTKQe9vdCo9bYT96jqA676U1m0Ctg3ckqn9sALE6MRpNl6wIAQGVz/D2AMSZMdmsMzeSH4I9zTqCE3QKYV4JJAEEAGg3mVauzkNqzizC/Dqe1/YfSsRMn0+GjuMvBBlplXnUIwC64JfNnwOYa3Z6uyjDH+gAdqHMjgvO30zIul7ffeQ+fu9PS8nJqCWrRrjGUHlFhVxWVv4ub5eLiUvorv/xXAb7q6Stf+gM2MNCFEhAcptgsDLIZWGOddp1z2GN8N/5Xi0ldDUaYwBETzTXETnJwCYo1xO9cjcv0s5husUTdsK4FIMUzAigx5ymLWU/7AGQE0RBWAGHhepmBsAygsVaFK2kG0SxXWQre5DWNMkIlbE/+RHP4XtRZHDPwZR4fd43M/TB/XMw9iXLiUrF0+MANKfrGucCRwJDnwjoeBagE+YpzMnE9A28iQ2PAqTFurrgEp7fPnEsvv34m3ff40+n4qbtoD33lWasVaN1jp1HcD3Fhfz1tEIS/wT0BUpm0bigwHFXS4cNH06lbT4UrozEijT2mu6rAKmH4IibdPl5qqGfqlmv5LgCdrsCyh3uycmmjqKT6KsDIq4foedEvfz+FG3CMpxo1lRtf7afAX7SJ/vuMn+t5+KKLZcgD+Xovg8mCahkwc5pyv3hQJXN8AMTGeO/q2jyZcd6ZjaMsMmKQseCjN7NsOLO0vDi+ePGiw3m9br+XqZRAKYE/vwRYkcpUSqCUQCmBUgKlBEoJlBJ4dyWg8WAqjt9b+43mWbZJgjql2Rh+hrt7Wxf29rYvtprNnm/uqzAQMCwmGKPs/NgTQeLcUrFBMAyHAFXBzvCSTAz+jYTTOK0BuRlD3+cKQyf4ClTcpGxjysjwas/10jIG18GjR9JXvvzV9PorrxGDbDt1mouYLtsYP4Bsc25IhhEGy8fA/DIaej1YA9i3Tc4nI2rEeJedBiUgG1kYPQJhNBojECOXc+PxaNAJ4MnEkUFRpwDkRQBnGst90vGt9Y2PHj986OriXPrCOnsKkBVAgQ6HM1VsG2e+Mr1nJKBGxthOW8w5SNbREydr84vLdTFSGDfgJY05MhxhB8lbYH8tsFsjRjSqAhTD3Q305ApwyjKuuE9z/hA61KaYF5kNr2Bws81jOsx1wLH6Ceo7aBnOHyz044Bh7mq5AgqwBFBWBVMAyRGcQLmq4HLo5NLSWjDF1mEFgVFFItp4xJBaaOfdWWVKLi+vpg6ukp25hQB5llcIoUe+InaTzJvNrfW0ceVi7E7Yg/21s8sOlOTpAbQJYtQA2OozC+nWU+9LD973IAH753HHnKV5zE3AGT+W49H1wV01ZbH1celrN6vpP/yP/na669bD6e/+1/9FgB4CG963DgP5j2fz8xPmOWH9AcoMxSaoAWDHXNYTzplkHS2AcKrhPuuGYJdzVKCFegVVfC4+nAfiIhDjvQCNAMbiHDEqUqapH1xZQ36WVVzzgucmd0v0CcsQRBfKYSWJeswfbbVeshf1mzd2kuTa9TaSJ1wKbTwpX8/PiBT5rPWof9fvmTFnD5AvmmQfKNe6jRHGQER+QSFlwwmPZA7GeCKer+wAPrv9tLezG7JngwlizM2kfhfWXwTXJw+sQ11qHdcGLyXaxCfrMYYQemNsZRPubG+mK9PNUYxPt7rvUOiHuwdXiIxXrzUBRhfT3NxcOnnyZDpx4kQ6f/FcevZrX01f/coXiSF5DtrWHq68BPKnXaEvxEZjl9Zol213s4a6MSMpj3B7dJWXLYyt/R3jxc+8AQTOgfrVJfVOeflptzOo6cgFCMq7FqFbn8EtMl6ImF+XYX9vyVzLssaveTwW+GYYqLmSZvl9dYhB6RETb5ux3aIk3sBU+ZXUaO/fv//Sxz72sa0zZ86k06dP23Z/N1htmUoJlBL4c0ogr15/zkLKx0sJlBIoJVBKoJRAKYFSAj+KBDDnMBx+8N/zU5ssipRf4Bs9PvPASofnIRH85Y88eudMvfL41vr6I/icLMs8wMAd88K9Ouz1qzMY1VhlGDYYbTASsB4CIIsg4Bo6GCkaixou2dADhOK7Brk2noBAsM1gnnmfjNwn3g1GjXHJ9h9Yg022GDFz+oBhI8C1FqCXHK4h7pdsFDBlhuH2MwMzzb+4MCw1Qo2VI4NNoE7mhddtB9YTRzcb4Dt1kjXcMa1XBgJss8poMGInAiWnORS7ni3Pzc9119bWXvz8H37tihHLMO1oiCha7grHMr1nJOCwOfJxDH3cf/hI7c67753pdvuY2xVYYvV5bGioMZWjZF5Bdyro5SbHXR7Dwq7Cs6myI17lfbiEPQZLaT/g2Bvc/2Pyv4U+L/C5BwP+fly5TpB/FZ1bpLwVpgmgWWUfM7PDdKr0+wAAgiAUADZbaeC+1nIHScAJd5KcAfgCuEu6P87Nr6Tl1QNpYWmVWGlH0z4YPEsr+wG0FmG8wBKbBSRjh0EZmTIznYN7e7u4Ue6GG6QgxSbxp5wjAY45B2FzrqwdTk88+XS6h10P19b24Z7mzo+whZiLDY4TgCyBilhN6IA4Af/BkHWtmwCqbKT9y/MAJF9Im1cvE3PMeVZJbQLlz+Ji2QTY6czQJuafjDHkESPgueWYLNN25Q/i4JorWLhHxnB5hWt+547z2Rno2hHXmOOxs4FlkCNiYl0vT/DFdch5z4f6dec0PqJl2I5YEyx5Wt71crkW7DSeoaJY06wvnqXNlpnbbK0uY5TLMdpkPk7ivr2Z9lE2IP/NFc+bJ4NtlBet907OHxnNbEPjoSwjAcO8AqE76E93aztdvngpvfn22XRpfTvd98TTae3IiTQYV/kAksEUHKAPBvHfAHQ9d/4MjLOdAM8cR5lzsVsleReWltKp226HLTbDGMNBQweUzyquuku47M4vLKXjJ06kg4cPpYNHcMU9fCSdOHVbBPfXfXMAjDyGjba4uIrLZpuYdwtpee0A7Rfo40UJOiMDUfdIWZHuVCnkR0dCRuptMPkUkWsxDxUfJWO+62s6Z46V5SrnAsj1UZP3TDwvwCVIFkDX9GUOmHNFsJoNYidbSLaLbtajjMmkzzzt0+dqpzNTPXfu3HWXS+spUymBUgL/5hLw780ylRIoJVBKoJRAKYFSAqUE3lUJaHL8KWlqZcC6wl6UvfHXP/nhpY9+8In7WpX0ZL0yurc1GR64cunCkcpwvP/KhfMRN4jYM2x+16rIWOltrPM2H6PXeEcATG1ctASxjPwi06Nge8gkMWXDWPYJscmmRihfxNiycQTwZQwgo9cAUaS1Q8cwxg5EsPDXX3olvfXa62m418MlrB/smN297QDTZJHt7GylhcZ8GEgaswMMrhYsCY1Vk5IgfliiLzSEDycaxZhPqU/eMKIA+oYjDCgkgxGFwYTLDQGoMAxvHfV79378I08f+sMvfvH07/zhtzHR3pGuxpLGW5neGxLIY5eNZsd/ed/B9MBDj9Vgn7SILcbukpUm47/ImO4jftJcdWzgu2TQ/T2ujevVhgb1KbT0BHpzpB4IbPputdJ8AbbPRe5Zxm0Y/Y+AetzL9w56ZCwyo+G3h6jVcNQHRIBN5VwgXldl3OT7BKCrQ5D7BRhhCzleFyC07sAj5lO7gzsyQEUP10gNeOPuqcOyudRfHI1xlxP8YWMLlLhRHQcQ0uvidvfW6+nalcupu7sZzzlSPRCeBk26977H0mOPP5mOAaYUsfosTxalzCvrktkGpJRqo1ra6e9EO5ozuE3G5oDj1MatsgGYIutM4IYQTmlze5RmAMjmYHF2ALbdZVPgA/ZlqnGUwjMBdHOOCpg5IuIOsspkcwpU0bGo3/boJiiQLXBk4vH4hnzjnK0QYv6HEzR0IDCYKLfAMm50q/YBNzawXoGYfM/qMthmme7YWJRtvpjjFiaYHvOdlkyf9bkiuRL4nKwm2wruyRXWHIE0W4zcvWI+gbIhAJD9zfHFrOcdtlvU73pK3hF6A7YTeXPb89rmmmng/h12Ar7CTsBDXia0AEe73S55bSvLGP96gGiunZvbW7AQ9wA+2UiB+I8j2GXB7A3dkak1TuvoyibxyQ4dORrgl27xDHow0ubYeRh2FW6WbLCyiBc6fRizdi8vrqQ777gLt9pO+tzn/yC9+MJpmMG8OGEsYOamAwdYy4/eCsNtKw14wTHghcvZt95M19YvR7tq6AxqBJgKWxl5Cp6pG74UUc9ZkAH4MlArO7I5bvN7QIZjHjcBXJ8rxkJWsKhjTd3lerjy0tZ4SYPoSYi30ka/wVJrJxDyZRq7y/W3cQntkmUB0Q0G/VEXl9Mev+vGzz333ESWWugCY5JTMfY0pEylBEoJ/JkkUAJkfyYxlZlKCZQSKCVQSqCUQCmBd1EC2mgVvKPwfUrpr33qmcP/1X/2tx7vbVz+6KC78ySA0F27u9uduZlG6m3v6gI5CcN80K/uAlLpRtOGGaALz+LKMvHD2IkSQ0twq8G1iYwyDEn5EDWMFGxDDLWpQctRdxoc1aK7GoTuOokLG3m0djKYxmNpbmY+HQbomoM9c/jw4fTKi6+kS+cvpC6BpjWOsCthOBCgnzKFrMJVp9oJME/j0o/l1MnIxgJhVIOHBftDY1W7ViCPjGH0mD8YZhAKlA8gGQwLAbTaURxG7/zsr3z6O//6C9++SF8wu3iETBpaHqIz5Y+fWAk4tqapcQsqQUD5peXq+5/6YG1ze6fFmBKPCCUhgDd5CcxfWUKrsK3rGxjQxhuDWThcIaD5LVx8AFW9g6Nwx2mM7FdhpBCPTLfKqsH3H8Kl9x6AjwPqH5SVPmpC/PNgY036PZx7BYEaDXCfNn6XtcriHMHs0fcZWGMtwGYBZ10tGwDQnuP4lQEmGmof9mDqDAGkhzsCIQItw2B+CQAM+102r5ChM0wXL55PO4Adu7CGBOZ8dszcmwXQeOiRJ9IHP/gM4MUR6mXXV1L0KGSV3SLjGmxMwTzBslqDtjhxaP8IGZp6zKmL586nM+cvM7kBZ1gLBDv2YAn5fYc1YxdAxDiBAeoBXtSRnO0rkuCeAJqgiMnvphg36otxs+1Mt2B5xd38w3s2OR+zfAKL4nqRLMdPlMPFKJejs7cA84u8ERsLYCvnz1et02dlVHk9XClvKMdcuf7pWhLAGBdd+Phe1MuXeJ5VhSaqkzlmlvf9uImB6Xp+c0XncpuViqBYkWzrCDl2Ab10ea0xJj5rPLLcftob1Loqu1b20IeL+SUFoJmbJczNdUKXBuiPY9ODcUiAej5X0hHi19XR2fk5XNxpr/fnAMZ0X3ftl+2rTgQTGLkYY3J+YTnde/8jjPcIAOztAOBG9L/ehBW5yAaSAGZNfjckwn7ddvud6eUXv5tePP3d1IWFOKCWPq6cDfRTXTE+mn0hQF8wGa1rwj6UgmXOK9XQ9VpdabXZQdn7cKFDdnA87b+goO0ka1zXvZ774WqpKPmAoY0OMd/v4nu8zeF+n3kMuU20dry+s703nJmZnTz22GOjL3zhC4j7Hb3lmTKVEigl8CNK4J0V7Ed8sMxeSqCUQCmBUgKlBEoJlBL4C5aA5lcgOlgGE8lUv/bpZ5b/47/57z9x4e03/1qzOvlwZTRc7ncHeDDCWJlhRzvcuvaIWTTG0NVNZ8iuZQuwXDTOic+VttevhaE1vzSPa85ympknPhIuXjVYDJk1kdkjMr00FH2TLzvAmDbG1NHY05AJvgUGkQayMckwWNIurIIW7jlrsBKanbm0giF/5o0302svvYhb1xYMFMxM+tCmLo2jYIIIzPGsRlRDIA4bCGIY5qCYCBsECJSFwajtynWMMQ2sYHHQRNkYxGKvDPq74BrZgqrXq2sYeY+cPH7La7ceXfjyq2c2NwQFprHIbD82VTbGs1H6jmH+Fzx+ZXH/BhIIfGE6PjGigAhLqwdqP/eRZ5owanCXlUhU1YOY0GONOUAHA+cTyLtK4KFKnzGFjMNGFfX6XeS7BzW5FV3GFbNxEb3baxIlH4bUEVhRx1Ggu7zfaLaX1CmMaVWDUwLY42aIX2YikF8aEGusCrjbJIYeN3FBXALIqAFUzUVsqDosGWNENWBgCe4KSEQMKvR5a2uLgPydOFbYpXAIYDwcUCtgSoDBgF17MMyuXbuS3n79tbRHMPYRgfmNZ1UHgDt87GR65P0fTPfc91A6dfIUO00CXPg0bTPGVAANADeeiyZnviRzhPmKk3XM4wHXRSgE406/ejp97v/+7bTFzoaGOhfk0XWuyzzewKVvBkBlCxdAISFZa5VxPXWZg02uC7YpIOswDmHRBxcp57PrQB467vEl2kQuQQoBHpNlyFQiQ9TByfV8dqGoo3jWY9R3PV8G0i0LlDTWgzyDeZgyTbbR52Sc+b04L8o0T1GP34sUTDJkBgaK/CmD/tgv+WSuNQV4lkEs6uGaXble7rQ9U1SfYu0rZbBm+anygsGXF8aWc5fKuMYzOwBksbMk9US9PCN7d2NjAwYZOwEzvvO4ss/gni77bAd9acD40zVWfXqb2FsPPvx49GkW8LYFY9C1WZkbgyxijHFuWwp2YAajWvzOWEp333Vv6NIFXqaou5VaK83OL6cFADnxMV+SbMBC1lt9/8Fj6Y3XXobpiK5uoqsBoOZydUG2XRKVmzDRKpyParmfA3RgnvIEwHxhMhzmcVd/BXAdI2Johq74ysPzGsCZCf0C42R22wFA8fFwfIJ13s03nLADPgzTpEtZO1zzN0atMzs/efLJD4z/+I//eMILJIvhWSHLqZL4rUylBEoJ/FAJlADZDxVRmaGUQCmBUgKlBEoJlBJ4lySgMeDHF/ARc+yDjz360HBn+y9VxqNn2GBvdQBjiixdjANQqnoboAknsmalCWNsMoMBggHnzpGCZcaWETxbv3I1vf3mm6l9+TLxjFb57A9Dqoq7TAMAAO5MGN0VzjE0MI4wrDCusBazQYjFpFGYYxphmGMECl6RE4NPw7SeOjBeZuZhKeAWtLCymr7zzW+kDZgOGoQDGGs9XM00nlpTw1HDU5ccWkBdGSSrYDhVCAKNWcQRY1rjjmt+cK/Tgor66Dq3arAMdPPRZXOyNBmNHsW15/VP/9IvvvA//r1/smE/SP6dpyEVVpIX+O6hTD9BEnhnSLDM0b6Z+YXaM7/wsfrG5hassDEjXZ8IHjHWM9jCq+4sSRwyxxZcrMpOltUFvt/KMN8Hi+YEOtkEHLuEbX0FlhebOkwONtu1eQCIU+jx3Vzv1A18X2sMdnd3ZaiAA+Mq1uzo+gYywkwDABsPaI9zwQ/gWBOgTJZZDaMeYxxAYTFAMV2a1WGRBVQydPXatWsBQNRnAZuYRw2aK1AgUDSCNSM4duH82QCSBwAo4gANXCBvv/O+9OBjT6aHYY8tr+IqR3wzQTGZODKEJES2AKoFoAJQ414PoFpAaRsWmIzKS1evpXMXL6SvMwdfOv1CunL+bfbzvMRMI8aYwARTt8+c6vWJjQWLbINYVzMwfHBHJT4a8QGrrCUB6AH3kDlAcVYk5BxaE/PR9aFI0j7pe8wtlwVc+oDWI3ZV4BtcI9C6N+KeYFKekhkwcY0wn897zB/AJds6na7FffOadE80FW2KE34UZZChuHT9mmUUiVpc3uKeAom2czPgRgXkf2AXXSsty2dFYVy3WFEiv9m8Hy3iuuuin1wW5+QT9Oqxg6QulcrN5LE4rwFM6ZpZY91TP7yuKybCi80dhsP8UiJkQv2yt/owDV1be7hCznUAaBsLUWaso5RtOX6ybADUAELthuPtOr5CDDP1R+CuD3vQ9grGzfH7wph06pm/P1rtQVo7cJwXK2tszHJLunvjSnr95RfTK7wA2ea7Lzlk93UBd9mHJc2O2K0VBpn1Nui7rr/qjlvHWoff7adjZ388H7BBgEfZzeYJl1MX9TzMlsXSPgIbqxEfEO7zcAh7rCZIFrtbMq8I3TZmi9nqNjEKR+1Wp/7oo4+Ov/SlL41xTRVgm45HiL78UUqglMCfQQL+ci1TKYFSAqUESgmUEiglUErgXZUAtlWkqf1X1K3V6S3jKmHkpLXOzNyHMOA+DLNqdaQhjKWD0VAfxXaQvN+HveJOkV7XmNTIqGOAzGPEG5y/y65pCxjaVzGYdd95+02CP1/bSvvW1gIkk01WBSzQ6Pe7BoXGiqwY6V+eyyLALsGuxaLkXNbIUDdNgQMMPDCIMB6tuyP4trCY6jDVvv21Z9PG1Sth0FWIvVPDCI8YZ6Op649tpiwNfS24hoH9KaMw7Cb0ow6DLYJ3264AxGSQDKvGeKI5kM+aY2zzNmS1O2BI3PmZT/3S4jeJr/PPf/85JBg4YyFqRVqmn1AJqEtCogtL++qf+PRnWjDHqhjL42aj1ccoJg4R6FS1uh/9OQxTS0DMOdJC5dfQk9vQmxPEUiIYvyb15ArAwwUM6W2mSo17sM4my+3ZOalYNdUtGF8orrG5ZMEI7DoXDWovTOKuqoJRQxQLYhbnBMFHVyO+EiASLl2hp+4WGGAEAJsKiRoHWLHbIBYSu0Puwf6ZncXtDZtf3e7D6Fq/uol726vp/NuvB4CtC5xuyvc/+Gh65uf/MrtV3skGGCsE6Cf2GTvNfumrX0vPPvv1dPXaJnMNBhl1gHUAeAzTLgCX59uwjmSQDQGie7BHjR/W7sBsI15ga34NAKMHkMweBiPKHO0x95mDCGIbkKTdbeKyR8zAYMgZw2mU2H6AcimYVI8tQuweABb9GPGpkEd3QdedWAeQWfwDgclQEfmZeRGzzHWDooyHpew9Nbm05CNPMNfz9zhQRgbgXH9iDYq1LS+OUbBl5azx07oiXyyf0zKmFRRlRFuDWSfDSzDOfD6IUli/jeN6oEjTZyMHfbUy63MMox70VabZ9PF4LJBHi/GhaRoBNOleuRe7RPZDbrqrbm0wljws6BbxH9GpAIwA1Po8o841Zewiz3n0p7cD44w1uld1bEdpHWbwHjHrVlePhZ64ZuJpH+trm3VWjEmgy/VW/RYcMx6eDF2KSfX9+/Ci7KX1y1diM4B59H+WuTDbmY/fC8E2Y8rJXhuNF5DXMADbYyfuSA8+vp7eev219M1v/DE7ap5nb8md1GW3TuU7gAFmP9hTOdWobzCgnTAz5xdmYzOIqJ9++XLE4P+2UXmO+f3iiNNsxmAUMf7MM6ZPvihhKvpvAUDuGH3d4+KAXWIntLPJub8cuoBle7Shwe/M+mOPPtH/+je+NgIAp8AodDoi5aGUQCmBHyaBEiD7YRIq75cSKCVQSqCUQCmBUgLvlgT8Sz5bhnzhBTzByNO9mJR3GFCZV+m7MEnYxWsAQ8YdIHNWtu3DPYyAzvHGHhaYBh33ahNi2BAfaX55QhyyhbTEDnivvng6XbhwKQ13uxHEf2XffgzrXqrDgmnymAYLJi/sB9yxKEOjewwYJeMAxg1NMbaR7BXyyhrR8NU+Ma9GpcH3CTC9uC+lO+5/OH3z2a8Qv2YLjA3XSUxCgzPXMUI1fMKgwiUUvxrqykGe3aEv8gA4aPRNrdgoO87DQCXgOegh/cVrCYyMZ6i+Q3OOw3w48syHPvzNfwFARms0YW+0V9+tcSzr+REkIMCCAghO1D716V+ub2xtV/uD/hhdxEY2HFh9gQBhhxnr29iE4hggBSpfWecj8HU7KMPdAGHsbDnZQ0dgjtXO1aqNazRhgnflHM912MBiHn3W529AuaK/+t3WOgC8rVnAMHQzGFmACbZF/Q99BawwqD0IAwwzdrREXdVbgRKLUSdl7ggKiPxoq/tdUEwGkfH3nI99WEQjmD8Ddqw8f+7t9Nabr6YuwAKtAHSbSY/Agd5x9QAAIABJREFUGnvyAx9O9957P6yx1dTqLKaz5y6lv/f3/+f09W+dTrs7zMdGK9pUh2k2VF50x70FmIK0ASYSLmz1BoxQPm0AMFinqUssqTaub82F/YBoW/RyN42qXB8Q+4m2umPhNiC6AeG3AHKauMuNgcdoGEAJjDP6Yn/sr8m+53kuezTHJPNeDmIvCGh/M/g0ESxRPvyLazwfQfc5WoafnPfmY573RZ6CkTU9txE+53Gaoj1csSyfvd5G7ud7uU1mn5LDon+2VUafzxlf0cU3zu0j64/lUDv3uYE8LFvAyTJD5h7J45oo61XvQDYRJj+sMl4gjMirq3sXFq+MLPQw1i2f3zZ2JM+yMW9ebxkH116BW/MBG4XcB7q6swzqviuGV29xh7HbwS23C2OwM2V89QHNBMVCH+lT6ONUSvYvPjRVgLOBvs4Qb2wyOpSuXrqaLkwuRJ9sly6abu4yB5a8TbwzCoq1X3fJHuBuXb2YWWCDgBPp7vsfSq++cjp97dkvp/Nvvh5x8PpDdzDmGXRP3Z5n84ouLDFTGzdLuscLnAyKec12hhz8vYM8dC2Fvxly5rY+xfl+rBGpQT9Waect0oI5oqhplY8sUfxBE36VFXaeHTRkxAGS9b74xS9OlCHpusrYT+VRplICpQS+vwRKgOz7y6W8WkqglEApgVICpQRKCfxblIDGd06aWloCOeXrGgriBcTWH4xmDEbv3/O4Wk0w0Iifz/t5jFwZXRpUJhlfWAlhtIfR5kWMFNkKvqmf30eMJYzgmZlOOkecsBe++Xy4am2t77EbJbFn1jCWCdysgVWHOdDswCarY1iFSyfto+x+j6heYguAc358wx8GF2CVhrnWp8H9q41qmq21ARzqqb2o4WRf2I2NQDMN4pUFC4b+VI39g1EUrB06Wwd86E9gEsAkG8HcEYSTVWYA7mBraKRSh0YrZl4YOQJ3tlFGD3bPPuR1il3iDuN5dG4L0ozSVZYkRTz9Guflj58UCTBw7c589dd+/d+r9YbAr1BkwBh0o0JzK20Cj+2nqbehFydh+sAeq66jD/4Nv4SuHwBSbnHtHIP7Bq6S5wFPrzLcgmVzKHFrhi0mWzMdgvqnediWGtmhcxrKwjcym1DkcFUkAFmwvAZOPoDj7iQDGeqZLmk7gBJV9N1zWTUyzBqwtIAzgu2Y4+dVUwuAZaSbJuCyGErs6DfcSa+/8h1A6m+kPVzUnNSt9nx64MFH0id+6TPp5K23wwjaB94yk149cz799//D/5S+/eWvMAmIgzaLWxz5jZHlvGvIeGMO4mEda0PA6sQRpPkoOUA0nXU3xRYxzbrjLgy1Q2kB8KZ/AYZZl+vk7Y26BFjnSL4dwJAGaN4ebDLnHBOTvgGyIVTXHwhlgDYGcBe6EUykAqAdNw3wqAQE5Jz/MlgB82N9AsNmbZiC9uakLuVfZXtewXXHQDaXwGIBWviMrFTzOjSuSTLRPDrzYxbTML7lei13ykDja+TzwSiPck3FxBcAEwzTNTDXR28olwpyPvoD2Bp1ez80xCqpP7t0Z7DQ9dAnzEtzo6xcB2umF/g49gNAJV1oBdbsp2uda7YMLWVUbzNg9td1k3bIUBQo6+FqqbslQHHkFTSzTzOsywK2ullubq7zTDQ7gC3bS3iueN78SktGln1mRxPASbTU75TThjU8B3i1tLxAzDOBMEBeqWX8vmjxssQ21nAnNs7eFdhq+CI7R6kMN3p1gHqXYJz9/B13pvc//ZH0/Ne/lr7yR19Av19MQ+bI9oTdOgW/YCvOuJ7T7yHgM7hhBOw3LmUBvNpf5ex4C8Q5twTNvR6/BAHJom9DRrlea7E4rCl68i8A5i1y7KI/F5ifm+z0usdzSHRSd3Oapz74gRExyQbbAIpCkY5RHvcst/JnKYFSAn9SAqxKZSolUEqglEApgVICpQRKCbzbEsiGW2G6Tc/4u0STcIJjlQZpWvv0xz/6+HKnfRf2i7YQkZcaBiqXmoEhrSFrTlgeGDfYX3HN2C+aAjLLdF2KfBhgGl9+72DYuCve+pXNdPniNQw1jEkMbd2zquAOtgVbiyPfMGx06dGoMK6QblcatgSFoiyYWzDGPGqUQwCK+ioSdbgeH4CsdXbpM9ZRi3rZGTAAsBoGmsV7bMh2wZiy6+BffMe047ssMdthCiOWB7R3BxieZsT1hmYBpFGx2TCeuFG71O0PL3zlueeuXN3Y7RWPc5snwz6iGr+W6SdGAlAQP/bxT1SXVteq65sbhKITjGDkCFyFXsw3Wu07AEkfACA+hP72ARN2GfhFlO999WYTl6vaLjHCnmu12s82aq1Xcb26yDzZrNdbbSbM8Xq9fQKVPUC8vXkYZcThBx3CAHcukBf9a6UmTMsG8wMgLQO4A/SehyIfBnob3c36juEOk4s2hR4b3F/dbDOfNPgFjIPdyXyIRCGCKYNhN129fD5951vPpotn32RO4SHKnLz9ffemT3zyV9LdMMcgucU8AtNL/+z/+d30r377dygCCI98wh0RI1AmDWkso4i2C+EEVON6YJB0JohAg/Mou2OSg/kJrg7w3WCzgVbqGwQel8smEfttm0wf9+ioUSbBngAzAFkANerWwT9ZRc7DiCPmuJg8p988Gin67rzyQx4BL+eZbY8UtwJuohyAE/4RWy6XSzmuL5HfZ6Kc6WPFOad53lKQ36flh/udjfOZG1JR1rR5N9wpyvmeIxlzG6bjNm2vpSrP6dLBQ0VRZnBThHwOfBXP2xRfBsgeGwGM7RLU3l1KrxKTTibVkHV2B9h+wG6+j3/ww2xyIvM34crILpesvxdwgzd+nSARQ0p17G4J4NSFiWbdewBVzo0BwOxxdrG87/77Q9YIJBoi0OZYyu51TJxLI8oNJh9y9ui6qtYI2u1QXh9XyzZ6r44vwDQW0BScqgZQmstxfa8DajW5506TjiubZqBn/F4BTDt67Hi6++570sGDh1QN2JGwJQHy3DTGFxz9Xl6z1UvZw/5z04I8pkpXvRUEzS71yjxAQeXKd3VmqheuD3ilVo1H2GTM2FMjxyTjnN1o0w6yYz2o4GU8pBuN2uHDhyrXrq7zO6jrKIecyh+lBEoJ/GAJ8JdlmUoJlBIoJVBKoJRAKYFSAj9eCUz/bOdQWKDRHuMvXcIGuIjbySFMhhq7uPGHPwZPE3qX1iGGhW6QMhI0IGS5aBiFaYVhotGhMeo9Y3q1cZ1pE7Os2cA7pTKTzrz2VrpygTgx/WuwTObT6hrG8Fiwymew3ASjPMXgkrWmAeN3XX5GgF5Y7uTDaNLABROLuE0aZHUCmrfn0iFi1mxjLJ197SUMKoJCyyKjlxVjO+GKo1Haw1BrYOxrvBiTR6BOw1tjyrbadg0m+0WY5umRXrGNIZQCDMLcP/J02MTgVuIx3frGW5dewHbdUooUY7H8z8k6y/STIgEN+0ronjv4gSdNGH9HFJVoECt/ZgE+2T6Arn0QmUREr0BNGhJv7BR6eDL0olp9GUv4OdC0FwDR8Pattfk+z/wwPvghDPqjAK4L6APluvuDKpwZOzJVoJiF0V9IhDzooBCC00uGEMxJdA8wLq4ZFF92TxNAwfrVJyBkHocdBLhlmpA3QBJAhYSL1xWAkldOfze98cpLnHfJUU0HDx9P/85nfy094G6EFWKDsRPtpN4BtL6afv/3P5eXAtonWCzIYBKcCLYUeUdV3D5hZAIfcIM5IvMGYNo5ETtaMjeNrWVsKpg1ADOD1Fk4nFoAIoNzOwRxg8EEY5NsADBDgJhu2m0zn2B3EfA8lhfgkbS3t8eGBHMB4IDvgJkzP7kemAznTifZY85P3aeV1cQJjLT5ER8ZWwGo0ZdIMLUEQAR0Yj7aPW/dMDUlrukGKgguW/aGW8gmz3mZcq4P01KjaM+vI3cOOuc3zXkzR7m+RMjVxmgLulFLzouS+Bz/XO9c17xe1ETtAdw4jl7PO1LaLMYAGRTsMfsoEDWAPWUZvmDQVV3Aa2d7My3sP5CaLQLdX15n7SYwPiCtmz70GYuIece4CVpdXV+nPcpQeQ1jvb9I/C/L1iXSlxdj5C310vFQ1iae4LubOsD8Ys32uuCXvy+2can1PNhigL5zgHWOneOYZSazDVYb4PEiZfiMSZdhRagLrv2TYSjYvLi8lh57/APpzjvvTm+++kp6w8/rr6ZN2j5G57sy37a7vJzB5ZjvHXaA7bOe2x5Bu0jIxzKtP3QewNmj88xEb8C+Ko3xcFInDp5KOkeLjuLSOaEcJFwBQK92Ub8+OVGdCS+UmrUHH354/N3vfmfkxhg3p1zuzdf+9LM/oU9/evbybimB95wESoDsPTdkZYNLCZQSKCVQSqCUwE+tBLQBb7QDexgOF/gT/gI7QS7xUnxmyPaRGgIYDOSDCyM7BOMrjFUelnEQQBJWkiwEXWtMXtO1yFONkRZg2Km778W+0EXz7XTu7EWCh8N42BrCBjgSsYjcebKFwSzLRBfHGtSEANsw0AQWbOpYQ7eCG5FAmfGbcMEUgag2MdA07qvNdASQrIeRfQ0GjS5g4Huxqx9WVRh0cAYy0EB769QRuB/1FcalRlq0HyMJThFWKGaQR39GwqAnxhORljCWqqfWVpZPPXD/qdlnv/FygGxkFL9TrmIBZfpJkwBjSTBwXCsDExovLy9PeoNhjehys4A9B2E1HQAgnsXNbY9NKXbRizl0YoVu9DDOv4nr5R+yy91LHIfE6FtEg/ajFkcALu7GfD/BnFlRXXQ5rPSGE8FdjXuD4MuRqnmcxhOT1aK7bncPIBal1p1MRpW6aApABX0UvDXOknPMTwB1AkMomqmFexoXIxD6YK+SNq5dSi+9+B0eAmRg6sqcfPKpp9Nd99zHNMEcEZTAdXpAwd/49gvEKMOQ55zMeR6p7oAvoh+2P9xCASoEZNyB02q9ltk2ul4iBUEzynPO6J7ZYHpcIbD7vpXDIGJX03DrbdwsAWVgAvXYkKNrvDXmsCB7E/ZQAxdLgYy6rpYwjWLdQFamIWCMQftBrOM8XBeVL30Jphm3lHmASraL+m/6zlPOa8aJHtInM5M8V7a57YI9WZ5xne8eTUVZPBHnxY8iX8x2Lgoq3VhGka842gUyFKfX816/cMMX21uUdWP9jr334khZbmAyQa6CZAJdypMe0S8BKoe6wu6Ru6m3vZ1avCTY3XPDEZ5neRKk8rPLvQ7ulLoi7nR3gsWXX34wFhXc0NGXbfJYZ5Esg2pCRgWTEBUNfVMu3vc5k8CarpUCvbrUF/cFy8wnOKf7rAH/CXppIbnd6EcVELYB03AwyGX5EsbfEe5+rHv96mobpuJ8OnHydvT+KoDv+XTpwvn09pk30zV26Bz2celElSuwy3xZMgTnGjmxSMZHu3EujVwUtNZRCq5DKM0xyWA18kCtDVNuGbdMNmqp1kbQNJvNVpe+tGnTJZ4iTmF1m/nZl9d59733NdfW1sbffv55O8R0UScRmHPsR0iFDvwIj5RZSwm8pySQZ/Z7qsllY0sJlBIoJVBKoJRAKYH3ugSynfeOYTbtD3/0azSGHa5d0PrMxz+yf21x4Sg7WB5mR8eZLoYVf6DDsoldHLFi4j/PwN7AONUdUvKGRngOnK0BAHOB/KZco4YeH+gg7dY8Bhy77W1jzGPw9HcBvXDwrBNDrIGrZA2AS4MvyosSaCL/W7hrhSvZFJnTjcdd0nowT/q4EO11BRU47uJqI8sBFzRAvjD0sLB41g/gm0YVDIJgyVgw/zWQNJJ1BzKfsjJvvq4hlq9hE3ErXIWGtXoVPEXcrTm/vLp6/hc+9vNfPXv2rfMvvfqWfc70tB/VEor+lj/+bUhAgzwnj5Xqo48/VT/94kvVl156cXRt49rgyJFbhjAeV3Dluh3wikD8tUVcvLogMD3cIvdjpB9oNtvnufa7AERfxb0SokzzVKPZvAvA63506hFYLfdgtx/ESJZWhfHeCqALoIJiAXIAmgyQTxnol25lqAn53MFSlzCbKJvROaaay2TR/UzQxbw+F/2Qxci5AFLElQL4lRHp/BszB65dvpC+9IXfS28RfwzELECkBx5+Iv3qr/2NtLyyxvwS9IJxRjlnL66nf/y//e/p0jlilFkp7aJw2oDJQpspNNhUssScy4LRASiZNyY3jfYeHffUtgqSBcuIMgQDR7FjoHN6gJslAJiuloAcTT23ecodN2NHWdpvv6rMQUEv+29/Zd8ZlN46nH9ea9FG52UAMDTBazK/BE14Mp51vL0fz1FWpOkx2hnP0COu+aygmd+jrNy5/Aw/zW/K9dBTT0OVpkeFEhdynuv5uGqybHN4DLFNC5j2yFXYB6OtAZ/Q10ium3z1hYH9iPcUlkN+Y4+NAEtRGkCgPmsfuzsCQm1vbbGbcDfWQ4YaEBRQjA0V9h06mu4AIJWNto37ZayfsHLd9TKAK0Ao2Y26QG5tb/C8wJvu7gCasrmQwZNPPpUWFxevt2P63oQ+5fYZ+8sXI0U7AZKDxba32wsGmaxFGXIwNNPsHK73sNcEd41XltlkyAnV0+UWZ82Qle6Vrs3uhGreJu2coZ1xjTng3GqiZzOdOTacWE5rBw7CTD6Yjhw9kQ4dPc6OlosIDB2lDOYr3WCuIG71KtqtoJGT/Qw9ju9TcFTEj4sC2RxV9JmglNUJGCjilSYLDNsKQFkDpvUO2rSBKy8OxiO0O7X2799fvf2OO8ZdNqnZYXMKpENlagKPlqmUQCmBkICYdJlKCZQSKCVQSqCUQCmBUgLvqgT8w//7JC9ySzMBUCtNtjc3N1+qHjn0EqyxB3FxWfYZDKURBl+F4M8GKsZQISA+b+G7OwBQGCgaaRqiAwI8AxxgHGFMkDQ2420/FkQVf8gKJkO9XU3L+w7i+nUljOEmbi81WGWXL+6lLdhkswtNdkprsBMmsXIG3TB+dJeyjZAFKAeDi/KscwCLqwe41iOm2S4gmTHQRhiCxjCam+ukVepZv3yWejSYjSWG+YL9b2Dm2BFTI4mmaqzZr8Ko9XvB4BHYG8BaoQUBBApCkDhoAmKMVyfNcb9/eDAar508cQv5vogcs/VTlOcDZfrxSgD9uckqZefKdMvJW2sAAmN0HrKXCoBHcb25AgC2QvwvqI7VETp80A+28ywW9RYA6yIMs9s5ngTAeYAxPkrPDpPnEDqzQIw893VwLnGoVSQfqjGyv9oa5miILmjOF+eHgG29Pkzugud57BagboMvo1txDTue52VbEeQel7gaN9VPgWAM8xDsBGZXE+BhE1bWlUsX09m3X6cRxpFi7gHMPf2hD6e1VXaQRWeNDabb5B6bYHzjm99O333hZcpwMsDWYu7QxFQFyMsSQ/MFShAANE3axE3B8GDDsHwATjg3+cF9zByK0W1PoER4g9wAE600u3wIdij9u8ycpuDKeId5CAQSYApssj13tsU9k77r+qcbHCsOGxGwrlC/c6lCmdH+YBPZd+Igxny0FllVHEixnnFdeeb7+bplTKdmZuZZppdI+V5+dnphei1nsMwij/ct1/K9nuu5+b55zH/jc36PZFkAgMU9y/IO7nlx2+emzYo8+aGbfzr+jnkV+emCOgDo8mXFgBcGbjhi2UX5gk8tGIxvvP5aAGhVVHueXU9l782wXu/btw8ALINk6qXtMdajyb4Vurq1sSnz8iaZmieekV3o+Ez1oqg75gLtchdT5wABvOgbMmNNFuBtwGjzeT8+Gy6Q5JCRRpQyxj/rujLRpZfWoKaZVahuOMFs75iyzAOrK+aFLvcz80u4+C6lhZXVtEassp3t9bS1sY6s2IyA3x39LvHVKHPiDrKKHqELulqe+ucumjLqjJkniI3rbxXgl9nTWELVd4JBOZmwZ3OaRW9lkm3yvcnYbPE8e1GMeb/U0wW78tRTT1Xefvvt9IUv/iFZrKxMpQRKCRQSKAGyQhLlsZRAKYFSAqUESgmUEvhxS4C/1MMqC6MeI2Hn5ZdffuGp++/+Tm9cvcYf+kdlEMBuMd4KbcVwwgBhH/swnnXh6e3KfMGFJ4wKjAsMDDxMwgifAFbJ6sKmwcjAtMHoasAAMEj53NxK2sIVKMcYmyMujqABRvv2ALeYrVS7sJHmlpoAZrhdYjiPdLuaA2CLv6Rkr8k8IegXBtsGcWaIo5x2MKwFyGZmYaPhEWMw5zCmMLTdIbMw3hS6xpqGWrBUNAhhrhg3p2o+M2B4arRlQ1NDmqsAFtkIxCiLoEeChxELaYk4PgeXlpba5Opi24kQ3mQIlSaRQv1xpnBuKxrgMA73HzhcPXnrqcrZs2fDZXduAT1szxk0rIUWzAJeddDdIcdVxn8furCGK+Eq7EF2rKyvAB7AFqvM4R6Gi9WYYPwwvRx8dMIU58TXEtTRwNal0Dhigg4BPGiMo1cCShrmgkMCCru7urLhRolrscm86qGAk3GZZKH1MPJl1FiHemqwewG13b3N9MLpb6Vr599GA3meOXfk8C0ENL+bXQEN/N9MA8DqXn+Szpw9n37v9/8/HEfJJ2hF22qz8xGQX5e3cHsT9BJs0SVNUIY5AtpCfYB91glZUkaa80OARzCtz26V7VniWgFaR8B+8oxnFgHIAdcHG2m8cwawkB01J5JwsryEiKxCt74MrkzSbGWW4PLuxshcpJ9IK1ztlJNguyw0n48yXMlEI8MVE6TMucp3WkT7edY+8DGmFo8E2M0BeWTZWoYpx9winycxafNzLGDxnG1xPJRJXjozQOMD1gUcGfX4uEkA1ASEEwAM3SAjsvJ52jUWUKJuGWLUENdtCblzHu5F3uI82uSJzF0BxuxyG8AiLFrBxRFyN8V6S33uKNImzuPrL7/EC4OraYadS1v0ocM6vES8MWWOm3G6Ruwu2X720f4qhdg5mIVW7qy651w5dstJVCHLwdhzjluFvri+KkddOk3qpN8HI3Sb0sbqfVwDHEYstdDforfqAWUqFvpF9bQf5KmF7tB2weAJIFiWBeVy37GjZTHf8GOOezPt2ZhH9TYbAaAn7qS8CEC2su9AxGBbZ4fMHUCyrU1cfgHIBMq6uAELlBm3LJhijINxAAXvbItj5Eg6J90lFKC61evtHWBTgTkYxFeZf1d4QTLD78gjgJFH0CH40ZM3kMWb48moy+hWcE+tHj16dPLRZz46+fIffXG8s7MVspqOrUIoRlbRRVKWxdgX18pjKYGfRgnEn3U/jR0r+1RKoJRAKYFSAqUESgm85yRQ/FFe4w9xzYD+t77z3avdT33iJZgdb9Gb+/q44mDaaBzxRzyGKkZLP5gr7bTLbmct3rCPYQgYL0wowHhKGUwj37iHLd0Jg0UWQzYC2cEP95i1Q7zR3zqLaw9A1wgDf5Jdz2bY9a7Wxc0Hhsnm1g7B/PcA1Si3U0+tbQIzL84HoNDQVa1C4PA+eTB4zhP4vzEzRx2wwSYLGE8TALZOtGVgHCaMPXAE2onRQ1t0z8FCCWPQ9haGr0cNE2/HNdyTdPfCx4Z+4GZKSZrdGHfBposA4ZPJbJPA7LAXjiCkNzDyhhqN0/R9jZ/iZnl81yXAeFSrAJxVfGMre3s7k0PHbsHIdtCq/UazvUd8IhECKV0LtA5soDLL/Fhm3BdqzdpttjgMVyZDMKoEN0BWOcWeHoMZ1AyRxGMZZPAoIhCgEzcEwbyWgTKU0gS4NAurpwfTRvfLRgPdphXqpvl1zSt0NIA0y5ExxFwUWCYX33swMc+ml196gQcpn0D8shyPnTiZDh08ErsG7nQpVyCDyaCP8KUr12gMWk1gdFCtNOY4hhUm8GEiACGzOrdXNz4KlB7HXOCHgMf0nn0Jt+roH2CgjDAAEHe4BURIGzCbDPDfmduXGsQQrADiyH4S1BNzUx4CMAEnOlFJytj+RdmwfGg0QfkFDQW6dDvN81YAI+JR2QaeMdkuk2VE7DJ6EeOQL1//LphpWd4zbzH/i2e9Hs9N799Yhvm5XJQYx3zt+sXi5vXyr1+YfjF/kYrvHr2az99pU3GuYgiO6U4rY8r112u6wes2qS4rAeBU6sUdFxkLhl28dCmdeeuNdOfKfhhdmYE3OzNmw4oOwOocLxs2w0VdUE921419nZubS5fZmfHKtY0Yd3VPuZkEaNU99dJUXFff3WDCTVGCKSjsxzXvu85bvkUUgJrf44UK00/gS9dbx6cB+83fO8YHUwZ5jAAXBU7JYxyy/D3HvVR3Z1tzoTtNGHIywWoc52CTzS6s4I7aTZvXrqS9nY109coFmGRzaRfAapf+V5h/A36vxQsS5NZXP5jT9pHfce5UqU7XqA+uc+rIaePavpnO7FH6BYg2lklWw810H/rZA9htcs3NW3psCjLmJUrlo8/8wvhf/O4/HwG0ZSRdhf4+KY/397lRXiol8FMmgRIg+ykb0LI7pQRKCZQSKCVQSuCnQAL+gW6Yn/TFr59O/+C3/snZX//lT39zMOjeTmyaE8Qjaxo8m7fmGiiRV5hI40U3H42GBkb2LAwU3+C3MbJbc8SIIQaT9ALMSNhcglK678Dmgt21enAJxsJWOvfGOkDYbsQQS9VlQK3FtH/lCG6TWwBxWzzLW/20h208TrjCpSsYNBrNxjiSLXHl2k66dPkaxttmOnX73enAoWMwyXppb0sDEgDPXfI08gUF6J/GWQUWgzFuTMaviS5hcGoYSp4QcBhiwOvCJW+Hbob7mkabhhiGaUWwwLICGCSAGoHVD2OmHcG0v4CZuK2U+J8tyB9gAEUDyh/vkgQY2EhYvaSZ2QW2m5uZtBhFxr/FLq144tY7AF31BkGSYEfOYtQfQMc7GMcN8kAOywa7xjJKw0fgFABF4xkdV48MGp91JAMHQa8RFDC2FnrID2oXrNXgzjooc9HzrIfop/AAIFnoqsBOgB3a0kB01BH5AESsxzhRw2EttdnNcmPjWvrWN/8YN7IrUUYwbHBvXF5aCeAajFeF50eei0tx1I5lAAAgAElEQVQry+goKgqwXJ1lDwJAlDHtrMFok9Xk89bhukBvyAN4JggiIGMC1IMhQz7bTpnM99w+qmFu6PYXbTYfc25nBChS7bBD5f40xl3PWGQUFvPNeqwjYpDxrGuKgFk1GETjcIsmQ8x9MB+eoe8w8iosMczwqG9C4H9B+Jh0gINOeAE4jw4X3Y6ZKDBTANhTiC/6aZtN3M4y9oRmZXfS6AlAXJaJZZivSDEmnBTu4JaVr2XAPV4OWC+yMEUdrC1VdxExxfqDfgEamt6JVebzjjmAIqMV4xFrEIwqBtQ4ZK6HAmOuWX5cq3VLtQ26187wGfWruFV20unvvpDuefBxxgZXVspx/VpaWuBFxW7a3J5NFy9epA1TV0b6el0v6asB9S9fvhyMM5pE+fAHGXt/Dwxpn58iOSfUN+eH1yXSuZ4OGTNdI5XjdRBOnZYfyREJAYyhawLKMWjquX1hnGF0ZT0RCDWn+peH1b4a26wAkpWz675zjrkdbGI3MGgYAgD9XV1dDUbZKvHKNpkvl86dxbV/Pm1vXA19llkW7DEBR9qRmWV5wxlBcd1TYUvXZnS5bjVPwcKDCNrivUv1eeSyTszCFnI5zvjMI5OzSOtaq1XvcY2dclvpAx/4wODZZ58db21tZIUoBDc9ql+FTn3PrfK0lMBPnQTyb8Kfum6VHSolUEqglEApgVICpQR+kiXwp/3BzT0tG2wKGBsYQr/7/37u/Cd/4ed/b7HRXB63Zj652esd1mDlD3ZenhMYv9era7Ts7m2DqmWDXYCszqdCPDDMKgwrDCMMf2PEyBjr81a+AuPLYPwtdksbYCgdvXU/dgOukRtd3ub307Vt4pJtTdKB+TV2JcPdTeMKdlmV3fW6vQ3c09oRQ2y4O0obm+sRD8eg/KP+VmrClli/8jY7sTXTAi5EfQykCXHSNHCJLBWGssaecojkfb56HtcweuybAIcGp8ZVuLiRz76EYRoGW7B6IMAMeCyXhWzarXrjILu0HaSKdm+Utqe6MK1selYeflwScBy0oDlWMdvrozpxmGCRVeqN1hpW9YF6rbUPtODWybh2L2N9gmur0EEW0ZmWu1GiJOIrUEmqBPNHp2LrxACVsclBCshB3tAJdeU6A0tkIG5mY10QdoCetafzRsO+gc4Zo0l9UkfVPegyARIIEjHx0N8MzBR6qPHsnBzjtihIPRhU08XzZ4kz9WqALbK2nKPzyyvp/gceoduwudBldVy3ziH3VlZW0q23n0rf+u5rlAOgBNsTGaQRH4EVgYEqrs+6WdMwpxK9BLjDvdE6ZRHZzmAwgZgIAspqUlYRPD76Tbv5pwveJmxUd7bsE/hvbf+RVN08w66CzjWahwjtu0BQyI8yPBYMMudgARjEvKUvLDORQhaWA3IWABWjUeR1LQJHyXPc9lCuMtcdFEiG9SibZkV+C7zxu+c+EwAXbbzxHuIxtz9ifDx63/w357MB3s1leSz6GPkB8dQur5kv6lOHKKfIG21G1mSi7b6YyHLK9QDYIPc+4yHwxw6sef2yPNqnfsnCmpmtpQsXLhF7DlkZ/wv2mQwv1q6IgSdwszgP8wr3XfVEPYxYZIjIwPu24epVGIeMZXY/zGt/0Wfb6tiE66g6E+cZdLSseh1Qj/XcDSVCz/l9IaB1vZ8Ac/E4MnSmKtlBFjKjKGAbc1ABIV9FxbVCRiF3ZW+tOYaYIQDoSLTbttsG+6ze9mG8OUfbgH4zs3O4/C/AaOZFC3NINtn6tctsILODczAbyQCWRfw0UGBBX+U0gB094fcE/ZipjGqHqXmOuTqijq1ardlFJnvKhftMLMU5GtIEhVIZDHZrc7MLlaeffjp97nOfG+FuOaJMMLhwGeb+gF+rQpB2RkUvUymBn24JTJfyn+5Olr0rJVBKoJRAKYFSAqUE3isS0IDxj/EwtWoYOLVuf9y988iht++/8646f9HfwR/ut2hsT4gG7Q5evFnHFpZdIKch/xnfgT2mu+UChoY7ToabjkYRTAANed2vzB35ZQO0MZRmYJ0RZ2xhFderRXYhm6tH/CJdXUZj3/YDrrX404l40bWmRllmCRh7qUFspzbAW7PdSLMdgoDzGRLUH4QuLeCGOUOQ/mB3UReGCWVhYmGIynYRbNAglyGjQSW+YYworC37iFFI33zIxto/8sjs4O70vEI8KULLcMvYZTCBsMLS+gunX37981/5xkvk2pqactn61mL7GU9TO/YGKSDfMACnQr7hzo/6tTCwf9Bz3Gc4pJf4aWCFNtKjH/wwTKalFXa1uw9k5+lqvf1htOxpsjwEe+sk2NkietICGMmPY8zLqhJVy+CYMwEooiFapJmusR+ulYAuGQCIanlOvXI3R0EB54zMmRYMxgAguO/1gYY7BrVgkvGP3NxCEIBi0T/1U8CCnSzJ78YYMmx8zjhPLZg5O5vX0rNf+WJ6+fTzlJVdxGTZfOjDH0sf/8Sn6CJGfbjeAcRMkaUJZcwur6avfut54onNOklSHcBgLHtN9iRlV2hnhbZPANjcybIiKxTARddL4z7JFKJzNNS5g2idNwIzXI/v9F2xeZ/Soi8VYo/tX0AGYJV4raWmLC/AH7aEjb7pWieLqEH9AhvRT+SWS4lDatM+1UfJK6a866wAiXPaD/3kvqxVM+ax4BuZzc+IcA+5ciYWYTk3JvNH4hBlCcBwwTHy3DLiE4PEOesHtbxz7Xp+rkWFGUxSNJ67LubM+YLri6PvuAZQNq3L+mJlDn3gQc5lDZpHQEWwVZf3vb1+2t7eCYaWbro0KJ5TpihpGrCIjuqddJWXC6fuepA1cjGqN35c9Azx6qLZxzV2awN3wy4u7jB2BShj91/a46YKbVhWjz/+BOOUY0a6bno9yxcJBUJGZpIMLJOyFWS277bHj7H6AjRjXLOs0UrGukH/lWPIku46XrLNYnzouzHM4q6AqXOCsl2/nSfOLR8I9llWl7jG48E+894QIFFZG1NNoEuX+w4vXmrMqRleyuACiavzPC9aDBXAaxf6T4F5fKlG1qdzVQ3SHZQxCECL4hrUK1tslWvEMEw9+jdg/WCDzWYdgBEMc7zTaDYGtNffo1XcP+v71/bX5wAl+T0ymZ2dqywuLVfvuuvu6vvuvLtqPY4BkuTzg5IdDc28OYOX/JSplMB7QALFH0rvgaaWTSwlUEqglEApgVICpQR+liTAn+HQY9yrLg3/0T/9v/p/6WMff67ZGn6p2e4cGfZ7x6qdat0A4rF73GQ44YidjPsKBrQG6zyGRRUGmUHEBaIMSK7xYxBodyfr7u2l2TmsJBkTjUlqE8WlNUdgcBhiO5s9Yr/4dp9dKfe6MMa22fEMRgHMB42pCq5iklPg/mDkNGClNcm3E7Y59h/GFQG8cd0E+8DAO5/WYJLNzi/iOsTuboaI5uEw8BlQja5gZPid9mmAalR5zX+eC+rp2qSRFAYq37mcn8PwAzDkUUxaA6FLwqhX13h8Ddyu2aWd2jS0Jp4q6vhZ0qXv7auyK1KWR3H25z/G+PzJYrQctbaBuKrQsQjqFfSaevX+p35u5fjJW49s7/bunVTqjwE8PQQ0cRJ78iCj1pAtVBdQEhyoE66MqF3oQwUQBHB4UhOYELSxH9jokfzuRx0SACtADoFirPsA10K/Qsey3qEcYaCLHGBDB+AhcOL8MqZTlC9pCGUSkBBH8pr9jfo497ubYly8dC69/MoLzDXAMRPl1Jkz73/qaeL3LQAKZGtZkEIgBu+wYNKcOnEs3X7q1nT6rSsAKMwtyqzafhtn25GDSSYoP+N7MMe4p9tzGgLAIARBmHEfVo0V2FCO/My2fYiA/gFMwI1JRCYEqOmm21ePMlnPpGoXBqiAC09McTDkKwCRWUz21VTIvHBzVJ6m+DkFuOMCPwS+7EIxDgGexIykLK5PdO9EJoJ4UbzXCrlO67N8r5mKe36PMskTYzDN632vF+Pj+ndzKoCgAijLAFbRN5QrsCXLKer0+Vi3GK+okzzKxIXQY1FnuFXKNEQS9kc5DXtAgICa6oGLIhoLG6uWvvvy6+k5di79xaPHwkXVPtoF12xj4Pls6DcX69zThdK6/XivDxAnq3GJlxAFiGsZ0T5bwHfXzgIcU3u9Ri3BZAvdo2zH1/LsQ5bBVLem/S9kcF0+lO13mWyqoWU6zwJbZUDzJgwZYCRrlJvl49ruOOaxabNr8hCdHQ3ZIIah5RVMktq1tLichp05YrARq2x2IS0sLQugZ7fLrY20fvVyvOQZM9fUYPmUyKnS56UMIOUYEJEhH67SJwGyeVD0NuvHq9S9i7zmue4vjD1kc4HfmcQpSwBgg7osztV9axU2eWksLy8Oz5w5M3jhhRedRgJvqvZ0hbFXPzwpo5CdaptF+sMfKnOUEvgxS6AEyH7MA1BWX0qglEApgVICpQR+NiWQjUkNlpvTTeee4DyY0uvr2+lv/Cd/6+Lf/2//u9/rtDor1YXxL+5ubx02vlilAr+rvzfhzXhtmZhh/lEuSIYFzBFWF14lDZgmGkBh1MCIISAxTANcbBKAGH8NNdzvkWObmDCEeUlLvLF397UhsXHGGDApzdGSHHtGgEvAYDyGtcI1ouFQVj9i4iwMCS69uZG2iaXTxXiTPTLCY7S/dw2GWT3NdTrE2qFMDC/MpjDqCnct2SWyI+KOIAaG5wRj6Z2EQQYbQwNLFgJfMIpgFGB6YJxpfuBlAzcDQlu92lxZWZpfgUwB140bWF8aOeYtjD2+l+m6BG7Su+tXv9+X60bf9OaN5wrY5BjelBjOUAbhk2pruO/YbekXfvFT6fgttx1tdWaf6HUHTwCYPlStNW7FE3it1qjNMM41A4HXYZXoHqwOY/hXBrjqathTHj+zGxiKiCGqDToFq2RYge4I3ti+2J2VY8QX41oNAMjknPCjTmRGo7qCme5Of8RYUjcFS5oATsEqcpMI8o6NidemLwJBMmfIFyxOyu4TP+r5b389nT9/BhAEw19WDu05duREuuXErfQH4IvmG5dJoICfAWTJ0FwGxP74R55Or/zWbwNIZzdK2waqCFsHN2PNc/Te/pii3e7uh3LXAcnctZYAY+QzXhgxymSvAZI7d+kMD1gxB9Aqmz4EAO8DiF/eq6Rjtdm0vKCHKwAgO1+2mDO6A7bbuIcyF2XrhDx5TmaRgEYwr8Ij3IlFuQDvxhQEpaN1gDvTNtZ5XjdCU6EvxTyM+czYmCwTcYRMzGeKPvJdoMjkdZFW63NXR5+P5LgAHMY4cq0AYXJ9tocURWagrag/6lEu1oq7osl7stDUsdwK9cuGeVSA1pWBMdmEcY3n1K8ebn/GILNcP7rHqlMuWpYvd3dUn0nnL22lty6sp3/wm/8oPYl7n+xcls0AE+EOhr6rKwJP6t8Ma7Nrou6FrnMyrkI21Ks8TFlC6lbubwbGWPjoS7D7aDdRvBg/ZkqMU5aFvY7xm/bLVwkmu6x86W2W81SMTmNTQG300YTEAvP2Udf9kJftoC5LCIZzFEtOrgno6YLboNNNXKxVzMqYFy3EJjOenfUKTivb2f5KWmIzg+PHb01XLl5Ily5dSBeYXzvbmzCf++x8uRvaVkdG6skQPRzgkil4CNjFTpYsJrXaAeR5AdlcoAF6VVfqrcaYF0bnuDfydw/gGgEPx/Vz587Vf/M3/yEer1LWQqx0CZ6zvz2yaOzy90mFgJSB/QII1fXay3/qc9+nqPJSKYEfkwS+93XCj6kZZbWlBEoJlBIoJVBKoJTAz5YEslHxQ/5qlmfip4bd11jf3ts799pr5z/0c0/PETPsEd6+7zNQMgb4LkHyK/Pzc7VZgC3fytcByDAMIJy0CIxPrDCYV7qgaI7vwSDb3dsl1ksn4og1MICNS1aVFYMxF7YWRou2dh0WWBP3y0odYxk6VsSdIQsv6OOjS1kYzjynq6WMCQ1qjRsD7w8A4rSfdJ/S9abtrpjk1YAjC+XBSMNw18XSZzX0ZXtwpoURhlZhaGqZaJdpNFqm57o3kabZscqJ30Z+kYBms916/WvPPfvla+u7F8kuLpAt9HfsSJ/9mU/K98+SbhyHPz0/gxl0p4oeVwyuFUBvqhDsCsJXa2Vf9T/9O//l/mMn73gYV8qP9vvjjwMsfAQXwwcZ4RWUoUld2N66PvGMT09jjKG/qEmt4rhrCBd6UPShaCPulehVBpHURY1fU0P3QxulzvFhL4BgRAqEhfsb98wvMqDLmC5r6lmwcJg76qnJeopyBTAsXxBDgGdj/XL6oy99Ll27hh0ueMIjwHzpwYceSR/8wNMBFOlapiscRXMPsAK916WtRRD8lbUD6SvPv5g297DNKVdX0grtDjdKvjNJEY1gGP2QKWZ7hCCiHtvHdRhwnjun6nzPhDMvcDtAHq31DB4KalVxr6yO++nkwVVYpz14PIDlYM4N5qqAoOuCMnPutXCjtq3KQvfSJtd1kRMAyXLlns8BogmWCLLFcPJMzOHps1QRAIlH15qcnPOCJ07l/N3rPlec+91PXKc/+ZwyIn8+FuCY42FO7ymPOOGHMqfFHDOg4a2cpt+QUQaUcvmCOVQEgIMG8gGpirFVP2yrbdAFD6A3QDJ32NVFUvdKQdtYe5HHhJcVu0j3areaTp+5ki4T6/Hyxna6/8EH0/ETt6BvrtDs1sizfrY3t9Cna7B5YfHC+O3CChwA+sjcCr1hDJ94/5MEuV+K+eCLh0I29tk54rl98TwS55zEWqpi+GLCW46tY6he209+Xn8mQN54PpcRbpQUlmXuXLDkLFe/FXXF/XzBn9eTpTiVBFxlK9YFkdUf67Zt6E+LTSqsx3nq7xjWc/LCKOMlUBsgeYadPHmCygBiGR9bHH2nAPJXiMU35vcLvR27c+USYNsC8hCJW2T+7KfrHdiqssc22WmUyTYBi6/NUEZzZnZ2cuLWk/1+rzcEQBs3iP3HSyC1ScW5rq3XO/SDvjhOWcV+UI7yeimBnzgJMKvKVEqglEApgVICpQRKCZQSeLcloNnm53uSlkO2Qa7fIJf0KD+Dty9cHPR73bnHHn34ccyfk6BAxGyZGczNzTbY1YxQRYBjGjoAYlotBD3HsPbPHXf66ge7QSPMN+1zC0sR66U1NysFK4wSbgGUYchhVmhcw+ShlQZZ1hDxpkwAPgGgZUNGwKsOOGbcGHezDBCNZw0crZElOKbpFEBYtA2DiKMx2jV8tLvCAPMcI0mpaFxrPIXJxf3cgyySDK5l402gJAAN82KHYrBrwfBotb68vPz6Jz/x8c8ThPn8159/WVNYgMziC6JFLrD8mXUOOb+TtAG5MGWSOEb59k2Z3sl+/RvPiU8yAIBbaApfA/0QvKylE/c9nP72f/53TjZas3+52x38KnbtxwkG9ADMjQPCMJjz8a9GYHO3cYVVRkkMZyCslICxbBKAkCkky1F7X+hXHSqAAAGkDGARJ0zgCn2MDzqW+8LcQG8bPuM8UYdD/wrXSYEPjW7AMcCsIg6Z88Pygv3Cc9Yty6WBkS+YJKPxlZdPpxe+8zXAEoKKo8fOQbxB02OPPZ4eeuhh5FghgHtmUQaQEzqfWWqCdAvL7G74xsX0yltnmFNtUWrmCQw2RW+cMT4CIQIHMsuiP7SFG9wWCFSSzDyHkOOEfgUxyr5737x+yMeXaLMSxNEtHVycTbPM7RpBz2eYt5ndg0yoKzOZAMBZY5zXtrXFnA850j4ZdIJmrge6jDrrI+aYDSQF8EG9Hk3KPVha3osPP2lSfI81w2ma88baw03XIjPFmDsY5LctohCQe3Jub07riDh1PmEWrnsrUqwXGQSyDPUnWK18z/nUK2oLAD4/FGui16hX0CMYgMYMUz+4PujDXEIv1Y0eGyD0YZLpzq7+uM6xkWK4s+6OG+mN9W567Twbm/BMBXmuHDiQHnjoUVYm9JoGufOlrL0tdhe9fOlKBKrXXdfdeq+7NU5jzT3y8MNp/8ED1DMFXGmL/fX5aPMNIF5Ii74HEEW3ZAv6EaBC5JkhiIBsg6kArASqcv8VLXrEuUfX8Zw8twzGn3GNecgNRyTmP22ieM+8eD2f670X/J1h/Z557hzLv3/4ncLLG4P3N1uEDgAY89OZm0/ziytplk+LoP6+EPK9CF0OvTLGmnHEZJK5FMGWhmc9ZorXWwCZ+5D60W6vv9AHhSQO2TbAW4/+oK71GdYRmci7AHR7Rw4fqc4vLFZnZzrj9915R/rMX/mr1dn5heprr76SBRTt/cE/6PZNyd9pyuF7Lt+UpzwpJfDjlkAxq3/c7SjrLyVQSqCUQCmBUgKlBEoJfF8J8Mc0JhfbQpIIe5/+6e/8y7c//alf/Pyh5ZVjw/7eKUKRzwKWabK53VZ1MCasN+CUgEQgQRirfeKIuWuehnpjBuYYMW5aBNJvYHTIHMOqSXiVhYGbmTkZGMPs9CLGESVpFJGngptZmDrSM7RRsQL8WoVl5q5oHWKfCRp0d4l5xvW+7Ac+wBnkl1GBgY1hJQgSFpEGPG2TxaMhLoCngSYrgAthkBZsINsWABzPaqjK7AnATIACcIz7xJ+REUFbJ6O5hc5M4+47bqe9v8OnTH+REkDEjH2UqM2HUqgggYlplRJmC/YXRvyEMQKZWfjwL31m5VO/8qtHt/cG79/pjj4GhvkkwNhcH3c09RLXMcIP4eCEITuuAm2McbBFsTTC1TGPAU7wXfey/gAdIdad17Q41QX1xdQQDOKoHgjEmEInpuc+EsaqnZjeEwzDzKbp1mUgfOL1wfLKYC4AhyxKcD7bUuiYoJHn6uVoDKgBw+eN115K7KAaYK9uzgLTM7NL6dDho7Ql9yFXKjghSIROU8ZEd+GJwGBKTzx8X/rDr34dUIyZQB4NfQGWG1gyUa/z0DIF5op+mn9M2wWrCnzHwP46pMoYmlRYSkTbEBdb9fGjlrrER9thDM5u9NmkYyHNsClHZYj7mmA4fba/ykGGmya+oJj1FTL1aDJPsJJsVywWACbem+aNTPxQZo6bo+SznhdlOJjcnV7LeePaTXmK53KJtsUyimTZxTWvF99tu+CNcgu2lYpDUg4ymIpYXTeW5ffrH8otvhe66Pm4n9eicGUEPdOFUZatCRXIdaEru+Nq2gEgO3PlQtqAbTZGz7owz9zlt8dg6WDOo5F0A15YWIi2Z08/ypn2SwN2QD1e171dtVdvCUUZz5ov8lo3V26UsddNXiv02GuexxjQltgo4UaZ5mKvP4f4Itn3IhV1FOfKXBAxypw+YPbr9ZBR92WLcv13XAT28jxnDiMv55U12DcFIzPStrZgP88vE5eMWGX79h9IVw8eZsfLM+kasckuXTibNmHd9bq7wsk8T9mMBW6vdHe4CFu15i7PlN1mng8BNieVxnCG+l4GPNvk91APd25IdOMOseBqx4/fkk783M+Nbr/9tuEXv/LVwec+/wdMmpxsa7TxBjkU9zzeKBO/B7h5Y4byeymBn0AJuL6UqZRAKYFSAqUESgmUEigl8JMhgXfsjRvbg/mgU09OO5N0/svPfuuf/c2//u/Ob1y58B9Mhr3lQW8He7SyC72shWFVizfpWLcYKbw5J0oYLLEBBlnP2DgYLp2FxQisr1FobCV3x5NFMIT1IEMlDJ+pwWSAcJ8JtgFbBuhiFIYkxjauKZggGt6aIVzH8KhVAN4woGVNaEDsEiemDaNCkExADEBPiwhmi2ibmAZGjMYPxzG9bGDMa1zJP8vGv8yIKRCCoaMBKSBgMdmYov2ADGMBE3JyNYGwUE9ENK9vbm7fKMvy+3UJZAM+n2qmkgyWbkKKkabHsP80YG8wBP06NXbD64z8Di1oD0BDWOz1dPCWW9OHPvqxpUcfe+rBzvzyUxcvX34E6OsuXAaPQN6Y6/cJIE7VYcTzuCcoMlkYfVlj6EDE36K8XJfFo7NWQ2w8cBuuE29IcIz2sLFr5BMsM1+OpYR+TF0sA5Ci4dkdkLrQMnXVh+2bei17xVSAQnGkfllYaGHonjtVBtBAfuPwOQfUwbdefz29/dYbadDr0n7mBm1Sh1dX1mD5HA4Y2z5nJbZWeh6iz3UHDsClu287lpZmG+kycxYPsWhfgFmISBB5LOoiAEVSLpbnHBKgcSfLCaCWLBr7bR+dL3nO8hzXZHsSCCuNA7hupCHlbtKuM9vDdHAJVmqzQ7uZY4Bpgj26UgtS6C7Z9ANQZr0y8IxDFvNVOAIhOScFH+2bU3zExhnwSaMPMkOLNsd4xhltpizlaTmCKiE47rnpRvQv8iGvqf6pcPG8fY+xK+5NdZR6zas8QjaxTuX1xfxZ43yU+jiPel0opymvcblduRzq417hUsnSxxi4Dmb3W0Eq47ypCwImdCPLDAEYj2wACLm7O0hXerX08oWr6dLWXqqxS+PuLgH2cam99/77WB930hyufLWC/ehayliGqzwyVY+MuWb5dCryGd9xY2NjKrfcftuEe2GWJ11VrsJM0UeuKzfnj7mDGWZpNPjG+4o1WIp8Mb/Aosl3IyEPzr3u95uSk9lkG/hYvimzSKlnml/Z+bzJEvL2KVxDbsE+cylgbvk7xD47jPQg/0MmbtrhnJuZIVbm4lLsdnno0CHcUa+m7Y114pOdTZcvnktXL1+SfQeTrGd8N3b4qIAVs0umc6hSneel0QPIqsEawzY11S4M7Oept0fz5pF3czAcDwHvxq+/eab5L//17/We/eofXeU3Mbtf0FA64GYKq6urk7fOvBm/F6Mz0av8w/mPpELH/A1ZplIC7wUJlADZe2GUyjaWEiglUEqglEApgZ9tCYTlw5/XuKBhx7Bl/f/yj3/ra7/0yV9cWZ5fvH174/Iv1XDTGfV7c/Vma4DRIh/CfJWewY75A90/zgMk4A/7+cXFVCeeiwCVQfAJjC7pgz/wyaVBE4aPNo4GpsAUBi6GCtYw3/ljH6NMo9sapiQJniEQP0wZ6/Iteb3eBjQaqZQAACAASURBVHDLbi8yITRcZjn2cImTNaDrZhhoGEL+syCNpOwah3FmHRiKfAtDM4Mkuol2w1jSuDLmk4CK37OBFSG2ZZGFUUj72beg3dTts0w3S0AA6mbjNst/ar/enHl6dnN+FACohY9YAiiOO1PWhrDGRERATxrLv/CpX1n9zF/97P7BuH5qe6f70M61rafgft2DK1hTwBPmGPjqGBxnUp+MY7BrBUjimGqwG/Tcev3uNZN5ZJeEEx/B5AcAO+qaO9hp+Bbt9Hjjd8swCeBYlnkFbARIZDnpouc8KFLkIa91uUGA26PK2KkScF+3Oosr2ikQg+sz7pUvsEnFtbhuO925kFmSTtx2ithi+2ALCUAzRzD6o1/OTfvHXBQc1pTGjw5wrJluO7o/XfruWeatjEsAOdtIpSEjQCrnqoCaQdsDBHKWF+336PwQUEGGsT6wsUaCBVdnF8WhQLkgloCVfVN+9OnC1rV0bmuQjhxYThXAOVmeVVh6gn3O9WIMlGUxJsV35YlU46MM/W5S3u/M03dAlRgbAYTpuJrXa36KbkQeb0yT59YjUGVSFibL8ON92xPrGNcdI5MukKYiT+gO15SXIIblRL3T/EW9riXmNUUcOvLGPeovnlEXTK59AS8zjoKZUR5t0t0dHCztwtq7wO7Ab1zcYKOSetrc2k13P/BA+vVf//V05MiBtL6+nmpL86nGeuUupzXW5Q47OUbZgGOWJ1i2RyyymBeCXLRjmxcQRRsLURb9tNsBnObuT/V7KmP7zvjTXOSSr4XsfGgqz6hcAdG36HdRQdwwW5ZNMQ4+X3zX1VKQ7HvnVO5PFrRPB7o+Lacoz7qiLI7FNZ8TLMsJyJWYmPa7Sky8hdZSml2YY6fLuTQ6eDAdPnw4fudcvnA+Xbh4vnKZwP6bW+uwmdmNNhGQv9oA64PjV63OAx7fC3uauIa4xvb6HZryGgzsLv0YwjBjqaxV9vZ644MHDw/vfN+do9OnTyOLMWMxW/27/83fTc9/59uT3/iN/3XS6+0Cv72j37YTqVJflhFfy1RK4D0hgRIge08MU9nIUgKlBEoJlBIoJfCzLoGp5RZmdGLXub30yV/97PP/5z/8jf9jeabT2dnuPxOGENjBgMj4uE02+IMfjxTdVCbwMCaEIoM5hoHVIIZLH0Mjx1+qhNGhIekf9wXAIFshm0UYx7IsMCAxRcLilHWm4ROMCQ0Z7ni3zpv5YGxocWkY8FyTTQNqBu/HGDfgdKVGS3gi4pJpOGukYz/oAmMyOHMY/P8/e28CZNlxnenlq3qv3qu1q3pHb+wGGjsBAgSxEgQBggRJcNNCiUOtHInawpYlOzwjTzjGsizNRIwnxhOjcYxG45Fsy+GwLNHDEGWJI4oixZFEElwAggSIfet97659ea+q/H0nb1YVQJBaTIIgcbP71r03b+bJkydP3rrnr5MnBXCw/sMEgi89Img0wAp50XPNOD3hrRLeBmHkgh/0NfRykTeYAXDpdSa2TgRt+gcFGSe9wo2VMDr1gghRKAwAAqSzlgAoI1VZLzT8GG6f4BDCqaGrETIHDNq2e1+67Q13XXz3W+69qT00euOJU6cvB4Dd1Vvp20zcrQk0bAA7NJaFaWTiLQM21Efw8QWBTZwX9TRyLBkinsfOjWZQRnBI7ylB2wZbuxK+KfRB3gWuBLKK51gY5vAm3xq+7vConW8sL8EA9dx6XmuIuxwxPFdC77JB26RPGRxzpSg7T6JzTZcRo99quNKz/2rVCh5aJ06eTEeP4D0GEKW3VYPlkgLFY+Nb0tWvvjZ2eaVKrgNf5dr2XVYcZ5bZtYgXDtKdbn3ttekvv/ho6m8TjByQbIVyeobFWECfVukQABxzyPaVT4ANAjZ0L8rxzKFxsAz0b74B410iucz84YKHzC+B6oGRiFF4+NxsumQCEL2fOIXIdJXlli4XbNkn6Min/VY2yk9wzmR7MT68Hzybr5xVq6hDmZCX5YIS9whR8CoDPOvggjiI9IxDV+pEG7Qdz+TFZqmbn9MPUhmTsrRPUJFCUS74UxAkPa8yCzZEhuPoA7JN+U3hGEKfB7bBf5I/cptxR2Z44EYT/EC2sBZphaWTglz4Q4J5rqQZYrw/ceRMmlxit1KWBf74T7033fv2t6Zz586mKd6NRIRPI8TbaiEzxyjGiT98jODty3aKCVem8N7LYf+JeYY+LrNbqQBZ9hC04egFY80Y0TWw0Ypv5VjxxUXx7IpMx7Cqp35leeSy0V8QLt/FMV+yMCiiUCzDSDpOIWfbyo2Ue3+PBPDsnKWMnmxRHuY8xx8+1BXus/5XA4DuBC3nJzTtu+Xb6Kvv//CkA8D1XZ+X+6JTvH9aLEn1d4W/58a3bI1dY/EgS6dOnUnHjx9NJ44eS+fOnm50uwsNYuaxupl3Tl9zmDl99WK3N8EGM5cxrz6Nd9kX0O2j6K9LLXvo8+xQe3j6siuuTlu372j6srr44otXnnzq2cYDD3wp/YN/8EuN3/7tf7967OjhIrg4Kw205fkifV6J+qaWwMtPAvlt+vLjq+aolkAtgVoCtQRqCdQSqCXwQglol2MqADBgn0wuLJ/5+X/wD//s3/2r/6nRN9Du9RZ7byQ8fbuNZQtQAE6GeQQKBuDUjysV4Y0wcond1NPowEA2TpFxvoqhIiDhtUYNF2FsR0BwYivpZZYN0WwMLVfxnrStjFejYd6Avkah3mWCCAYHJxtnIow+nLhGoTs3MxsGpUu8gg+NbfoTPGDdeuc6PZd19jQw8TTr4QWnoR28wVdsHADkl4Eyl8StG+w0DEMCIBEbpkWZUdbXaDXCvh2M5rh9ZSdll5OQgteISOPYwdiQsm6sAQI4Wrn+kQqrbnvYn7co1clmaHz7j3zgJy+6+ZbX72PYrp6aX75pefbC65bTwK4ecZFc+iiwQQOshgw9E0HpX+65aCt7/Amo2J5J/hxzdU7D2eQzH3uv/kRZwSmXtaGjAlgBxFBHUCwb3DAnMEQyrpgp32dASns/01XvoRttCuygKKUt8gRie2zEqSEvOMsmeeg8+oncZE8I+rlnn0zTM+fRYb3jVmLDipHR8XTZZVdxXJH5idmb+ycvpb9BnzkluNZe7iCl5fS6a69O4yOdhL8QgIBgoRME4VcgRVw7YI5ZACIKGBkBSMubsjOFlxjCj1uyKBFePZLRy6yf5WrKWw+yRv9QOs1SP73IJraP4TM3T2noApAIZvFuQU1yXDbpC04oswDGYnwkSpvKrhrLMiYxeDyLe9oyCeqZpFVkEedMZu1ZXPBD3rNO5LP50it6m+syJtDLYsrtWM56/F8b7/U5sN7+Wl7hR/1izHJd6+drp4yeY8aGU9dEAcWQfA9Kw/IIFrnwLmJZ+oUzF9LjR06D6A6le9/0pvTeH3x/2gQI2VuYT8t4Hhp83/fczMxMGhlioxP6FB690JE+Gkme2yi4BL0V3rqK1/4uzM8GYOS1QKvtE5Q+ziGEqu/KwOeOl0tXSxvmmwQ7pZHlm8dF4Dg/87wu85IXXoiVrKLPlpKxklfdR155ZmVStB9KGMVzvfwoeIh+q9fQkpsI/s+FuyP3xVxZ3xRB/1M3gYldahmLAf4IFH9UYb52OkNpbNM2wLKD/JFmMh07fqTv2LFD6ejhQ6vzs3PLzD3/kDKMB+qlNMP7amWiv7kyipye4PfoHOcLeJAe948tY5sm3PxliTE4PzI4NHvy5MnVd9z7Ln7Hpcbp04yvQsoJBXh+8sHXZD6/SH1XS+BlIYEaIHtZDEPNRC2BWgK1BGoJ1BKoJfANJSB4oR2RvX6w/zDOcBB4+NDxIx/4z37hY//zP/vV2ZFme7q3vHAvRuQgscB0LZnFy2oAcAzbwnhNAgTZ4MCaCMPP73nMHsCLDJRpD4VNpM3JdRiMtKknhl457Cmo7YMhrWeAhqB8YcBID+NLQI1aXGsomY8xQwu9psDZIBsEkEdb0taDLZINkgHpMIZ8Zhs+1jOGhrjPngqWl57LJoM32op2MCgx+rTgqG2fiINGYDWM2E3nz5/fROYFMmF4zb+DrFeyvRL6FOJ3vIokKtu2ukfSGuqOcdY/R5rRQswE4Teg/Pa9+9Pb3/U9+9967/e+7fyFmTvOXbhwMWO+ZbW/OQ4wO65BrqHLEsrKAGYtJeDTMmuaBFCIzhTjqP5oCGtIZ8NZUA19c5BC4Rg6rhvGlnOsiTsmnSbLrAYYaw1++WRXuuhT1g3qihlhPKs15glEZWPd4V+PnxUdFgQi1+fqsSX62WdA3qw30F4hkDq6jSxYmxWAkbtUsuldOnn8ufTM04+xhGuOWoJjQ2lwaCzt2LknXX/DjYAe7BSLHsccgb4itf+CL7YnKOx8CM9IwJLUN5cu3jeabr/5uvTRv3oQRoboO2Xw0jSYe3iKwSwwMnORDsq4Z8rEM24h7M9IxgZ0fjl38H7xZ+T3AbYYI2yAJde9BcAe5mhvdTQdOj+bdm5h90DjAa6yGyPLPgfaGaR2gwRBFvl2Sa2HoGPwoXbQj5Ahz10m7TjGmMIO3QxgSU5MysNnCiSAkNC36FjmT9nQljSkKdvqnxfRvt5N5kmbH+RmfaGEIJnJ/DVAyNcDqeha8RQzW17yu0c94BpZGkvNeFkmtNhCUVfwRb32bJ/c7dL76AtlY5zRjTmAnOfOTqZHjp5Ko9v3pL//Qx9I17zmteHpODc/E+Vw+AVoy4H252fm0+Io14ikRUD6ZeLs+Q4NjzDoLtHOPDqOh9Mar6dOncrLP2WSZNsBRsfviiwDBVT67PMQIWVtx+QSY3vNKeRbPMyyrHMZqzn7Yz7G+HFNeVswbloAiXFHXtDL9TaOa5N82xdQzXQyf75nfFeU5LMYqjLu8sZ1LIWmUIc/+DgH87zPuiBdgfhIwasTnw7G3PJdMcDulyNpx55d6aq5q9PZc6fT4aefbjz2+KOr09PTjQ70mDvD6NtrllcaW1nyfAQRniAG33NsEnOk2epM0y8mbDqzuNR7cmHh3OLw2Gjvi1/6YvrIhz8EE+v8ZybWf1ajsJ5RX9USeBlLIH5lvoz5q1mrJVBLoJZALYFaArUEXoESCGNwY7+zXUdOuYjFP5ojq+enZ6cee/iho2+6+645MINR1o3sx1ATWxjAEKFCn38lB7No4U0WlgP1sgGiMa0XgIaRqY/1WMVI1LCI5VvWiTIUCquFglyG9wf3YZjCiDQ0fKxjeUxJKcZZI1fEyzoNDD4NGY3JyKdiE08xAzIHH9Q1iLpggYaqjRmfybhJpjBEBegonA22DDIQ1wmnuABYsIWMGZUmmwOtrz53+Ogzf/Kpz05jS0Og6uhaRyz2Sk5fz3TLljOGqgJD2A7WwHJfa4ChIyhVf3vLD/3Uzx34yZ/9+deMb991z6nTF95NmJ63giXsIX7SBN5cg4sse1zuri6x3M1BRNUYAbQAmgy9qGgeS/VEXYglwoxP6JM6RFrXEb0CAarUL8oGTMdYhyEtdAGYoYEc9xjSAjPSKRtFaLDreaLBb33YiXPWIZiCLkXIyx5R5qu7YehDr1cBIi57E0pQHC08utQ38DN2rnw8PfrYVwBMBO7wZCHIvQG89+zeTwD2a9PmzRPUoh56K9AsH7YhPW1454xN8kjWWCIGCEVssMHRzelTf/XZtNw/SC8BinjMotSgYQX5WBtB6ZonIdvymquSvHO+h4yc0wyBu9gah0qPI0e6D/6Wu3iNAYptIabT2EAjDYKrD/Au6NDRAfo8gBztS4wHAJseTfLi2JiyLCs+YM53QiTpUy4vfzTHcXJuA5hU4y1vmX9lUT2npHlxT3/juaiU+QivlPf8wiPKkO+7LGg7pgq5HEGFH9zH+8pH/PO/SS8xywuOuXzXfOPH+QeFAH6lQ2aRq+PpHgxLOK3OsJTymZMX2Bl0Pl1xw23p+9//I+mSgwdzHDv620T+6ssccbFm2WVY3l0Sr1feIEst5akLGDZ5YTIdPnIUTzG8zWyXd6FgkuWJ55dGWVZ42+13hP7jkZn5rviPfsph8In8K/kp7pBVpYexH0bUXC8TtyE7CShDDpN1Q+/W9a0sz5ambZT2lI1HxPoLr0YJ+DrgpySrs/IsqcSP60cO6hIjHHoi7Y2JX2drbdmeYGdQjL6v64u3xvgL/iGh/g0A8o5PTDR2793TILi/2rSC9x7OfOw4S+J34jaq7eWvS1upMgH/2/mdtBseLmK+DLMMliL9q+Q1Op1236sOHGicOHZ8dXFhEVLyWTGRb7jP6YV9KPn1uZbAy0kCtQfZy2k0al5qCdQSqCVQS6CWwCtUAuXTPz6rkUExMPygjuvyIBsXcccPF31hdqTVzz/+7IVf+pVf+6t/9o9/ycjDfKh334lxgQmGLwAhnrBCWxhjxIvG80pjif+uldMYFFgwxce7eJrGBiZDNtorgycMUg2fKEoZjVEMFAwPPXf8w7qWU/CKLUKz3PEvmqqW0JHXxuAxmL+GnkvjLGDMnQAtADUAYMLQ0XgagHsNwRyoXZYNopw93bTX9OqRjhigBhaeRcaLwea2D9w32WovsUnc1u3jnI9LgH6ZKLBuxXBdp68rAQbIiP6Odl+nt23XvvS+H/rx9pvf+q47pubm3/bo449dTdyw3cTa2gYo1jS4+DLBwbp4uuhixfjgyKMOhX7pv6fsGS8AGfTDFEvHGD/BKGMNAVWFp4g6UZ7pRZPLmpfrOc79LHUcaLB8GGBCPdb4NR7ZxmSMqBb6q765xFidU3f1yhE40fPJa+na1XzkNtQx6VrPFcuJGHr9epeh1/0sn9ODrLc4lZ56+gnKqZtZLwWNOu2htH379thhL+JUUZZOR9vAhOg2sw8dJ/YRyyKd5/IDaAi/9scNRW+8anu6dNfW9NDxOfo6xGTXe8hJCC+U1xssGrVhkp5vMQedqOQ5Z/I7JAM9AlLKmc5GeedZhi3pO3WUXx/g3szqYjpELLKdg4OJtWZ5D0rKFvqCjYIXlrepuIZ52wLXDrBMuSq77MnlwDNP4V3wO7OXy/seMikeRjT4zzwLWtmN/JwXEoWUE7TwJDRVVSnjvXJZT1GOsY58ymdwLnus+d5QjPIhjdJe1Cavh/zjoeegkN9tAWjSZ//QIGVp24737qTKrod4+K2m83O9dOQ8QOPotvSWu15PMP4bUpvltl3oqXa+s5bRNfVEfXdpOntWpGHez5EsB0AkuGhMRt+ZjpObLQzQljsC266HQftj8wjKmqLfnpU942xfX5hChdAzpLI2ZkpfOaB58e7ntC5RBQXjalToj+93ymZQinJg5tYNuUqHPgYflglCtBW/W5Q1faJt9Tw2W3Bc+W+KOU8dW87zMb87HCTp5TLwSN9wuos2gdGCXz07S1+jLnQDjFbXoWl9ZZoVHt2C3ACennv2X0JcsW3pyquuaNx///3pyHOHkLm/l1psJtK4aCB2emntoO0pSE5z3sZy5wl+n26Dy2db7c6J7Tt2Tv7EB39mkmWWc7//od9Li3OzdCGW9styZtyLqg9m1qmWwMtVAvlN8nLlruarlkAtgVoCtQRqCdQSeEVIoLIP/q59DevwxOnzM089/tVTb3nzm6d1puLYgTfCENYDQYnc4p7P/T43CswgUok/pjHhh3s5CyRkW14jMRsjLrnRCyCWHVWGmOVNxbjMQBnmkEZRHNDleVgHAhLQWCXklN4HYZ3GE42jYJ87AQ8xreyNEgCGBgXPpa0xDgMYL4AvsGYg9Gxv2EIYg1qzNB0EWVLTnGel6aGnnzv8zP/7p586yUO28YuUGa9Yq/JeUSfHp6SN1zkvxMMPBiqizbN5at9Ab9O2XQP/9rf+j71bd+5765PPHvneM5PT78Qp7ApM43EwgQG8WZZWeqvEE9ffptHA4wYVaeoxJnYJToL6lXYDncg8OHry4J1ghbooCCU45fjqLaZnk2CsBm6LfPNMjrTlXQbnWS+fAGXQ1dBn6HoOT5TqLPhrjDrVsDzzuTwUz7PsgBlwAHQNsg7IQJsa4DZtjC95GMDoP37sUHrg/s9QZj6DZwAAQyPjLLEcTtdd99q086KLAlzI/bG3uZ8a7wLAaHH00x7Jh8llpAOAJ0Od/tQeHE+f+PQXcNobhEeAQjot+GR/7UTMp6ilLJSl0od3aMdE4afitq/KKQoFOJnbXQXMzHMzoBGuAQSR88LcZNq/bVPqgNSNtfGYYzlnmzFwKajlQ17IUcAjxgj6RZ4xno4ph8nnkQcwiJSrvDyvSxkYIz8DGet5UTQATGUTfZZeoV3OVb0oHavgchvSlBavjbWkfoT6Iaxoh2ZtORATyvq8tKMM4x4Fd1MD66kDMW4Q9X3ovWWWuJ8jGP+52V46Cjg2vutAuvXud6Qdew8QeowlstB2XEOXbRuZsIdrmpqZBvAKtCd0uwX4qJeeE8JZcZIllIcPH0p6N6mfbk6SAeEMjrYAze66+814pLUAynLsuQDy6FLph90rMjUvzx/OtqB8bItzKfPCMw9ibOWp0LLPjoP0sv5U8sxFXvBTXfN5BQDHUEcHo1zcIg8HYiMfjmK+z7rlNWSCTm5feNHfG3n+5ueZD68pGfQF5KxkE0GPhqzvrxQHFd1qbNo01rd7957G+PjEytz8/PLiIt5g7G0zPDLSRq+HkNlQqzUwhk6M87twC7+TRpsi505kwGpjfW7ZurV91VVXNb74uc+LSpbJJg/rzHhXp1oCL2MJ1ADZy3hwatZqCdQSqCVQS6CWwHetBL7mczlMAbrrF/s3SqWcBKKsF/pJxM2RU+cXH3r4oWN333Hnk3zkzPHRfhHm4ASGkz5ehA6PD/U+l+ZoWGss+Jd8l22FMYXnlYkv/jhrY2iUhSGBFaUBTE4YKRoqAg1RGiNDbwdpYp7E2ZY0IF3CFZiVFQQuIBrxikQ3fAYFthSIc26WHMpE3LEw4aIJnmvQaWhhjHarOD2AJdjrVSkao7PwQROxpG4Rl7ljx0+fefoPPvqJw5hzrh1TAkWIuZOQfyWmMBRDziEGh4GkaExhSqIgOim20oFXv7bvf/yX/+amZ48c/8Dk9NyP9hqNG4jDM6HTlLrhEkTijDHcKAnyjRNWsykb5IIo6gekadNB8KdGaigTD0K3ivUbT3OcuqJX6prAjca83Fnef2Zk4CfzITgQdKHPEqkMqNGmHpGwgDGNbqDTAkl6tejRZAwl6QRNdRgdC1An6GeVUUedCMsCSuohcbmahGL76sMPpmcJ0C9PAyyLHB7dxNMmgcE3E2/q+jSxeTNgLRg1z8OWDh1eVz3bND+8t2hPsEFaYmUt4gZeceW29Ln7H2OXzNOp2RnFASYvR475qiyVYfRH4TIBQr5c5gWZnHiuPDnpxBOgBjzEOIS8eRzDDspJnCbbVS7Li/NpYqiVdmwaTkP97Bi4DL4MMOimGGVMBP0ADYKU/bDtkCHjZJMx18krLMV4yQ1joTwyWF6Vy0wEjdIHzwJjyqck87yLnAqkUWbryfbKPWcaWrtXWaEVamiFqv++7xxziYb3Ho9iI5Iowtj4XvT1QnuWiyWW6jzv0SX0YgEPrwvz3XRqajGdX2ykg9ffml77+rvT4PjW1E+8xBYbRATAq64pJ9uFnmDXPMsrlxYBvciyry6xHECu7WrpqsHfjxw5khYI5u9yVPZfic0BMihFPEa8/G695TaWEOdNKBzuzCcEKzmU/ue5SPt01HHyuRDtxhTjV8aSR5ZWvCFiaLtzZMydEHG1tDauBR59+ytGQSqpVrKv5B48+zxkDQ/oASWCtnIxhR7RTryq154HsciUrmVCL6Br32KZrjzLm3QUJkmvu+IdmjOUCXK2LPWk47vLMv6+GQCE3rp166qg9uimscbC4lJjfmkRte1rDQ8PgVsODOL1NzLQHBhrtthxAQCNZytuoMEfd9pwMzo2Otq88667Fr785S8v6ekXDYa2Bwf1j1oCL3sJ8PauUy2BWgK1BGoJ1BKoJVBL4CWWQPW9v95qyXi+sbL+vFyVct57HeW1Nf0E97tm9fjpc3NPPPLVw3e/+e5jxLDhD94rE+wwuYnirC/DRGE9pItbMJJcbBYG+bLGHkZFGEIYDRo4GlkaEBrumBJx1lwyFUPLa4EPDUaNH40On3kO/ipDxTwKRH4saYOu8Y8sYxtNPMfKcq0AC+iMxnUYMpkS93oI6cFjnzXxPMdf/wEt2GmTpaWAeTxdbUgb7rvsdnjm1NnzT3/4j/70Kcy3mbC6sI+oaArh5cv6JxJg0ESKGBDdiBotzNRmc98V1+78R7/8T247eXbyBxZ6vR/Ef+/gUnd5ECAK1KBvAVvXwW3gSaNcdVF0VZ165pLXGN+iF4JOa/pBawKokSrdiGdSE8kiGddqLbYVbGVAC7CNfwJbEAudsp3i2eO17XlEGbrlUjaqE9er6FuObxTeaJWuqsca3blePgvkeK+qaNQT3y/aBB3jjCdRbz795V/+eZqdmcJA1svNw7he7bR7736WbV2V2kODma4MYIQ7l6Rnsr8eeKtg5Dvn6Lv957mgzGAAa610xVWvTg8++OV0+twFNroYtNtRXoAhL7NEXrAZ8g0iECIF/7Ybc5j24N+4VwFQQ0SgK+aRI8/YCC5aXDCn6ZK1uZm0lxXKE028ypYXIo8tP9CKvMTSuauMPZfDdu2dcisAmX30eZYl7FDC+5wsty4Ty4QehNxzCemtl1dumb4jY74AifUK/VK/5HkfqaonXyZ32wXugpt8n99B+d3nc3VK2fl+k4bLaEPPuHdZY4+8he5qOj05m05NAyAObk433HFP2nPw1Wm1xbizQyhAyhpIk2XgOGQQdx5gDBAmPMgWAdkG2k3G3E0QjHGnjJtpamqKDSCeTgSShyP7yDJiwNkefyTw3liNd7/5ngDIXOKZ+czjX+RgX0xFHupXSZYp3o3qv0k+Y3Uq15lGrpvHiUz1RXlDJsCukKdS5IG/RJyhSoUb6QAAIABJREFUzCfrmiKfcwCd1ThZfyN/+TrriLNkjdeqfEUon6I9LqN92qXNrAeZ9xJTzdalEwz7M9iRzzzvShv+8pTVDOL3NQbanT68wRpbt++I31PsqIwf5Wp/u9XGYW+gzbzqoBZt3lMDeK91qN6BBcg1Fmdm5xaRY99tt93Wf9999zXwPESJQlJwEGmdoZJTn2sJvIwkkN8CLyOGalZqCdQSqCVQS6CWQC2BV6IE/HKPr/e/pvOlXDk/r3iDD3U3nExHTp9LDz305dPvfOu9T/DhPrXU623HitgbMb20gi24orWeTcNsMGTjKgwVeAnjGxgtgwYYPAEWZKPWv8xjDsSheanNTwkzszHEo0xHgwcjOowmnmokaxhr2FsDzwrBEJe0NdgJr5+lRXpCFMNFYzC8LcLQwqiRdQxarRltapcjabRKS6ylCspOE9AZaInaXThy4sxTf/DHH3+UmlOVtMr3X7YinyfC75wbZeQue99Qb2KcNvYpj1Gpk0ewPHeQRKawBcXJ8IK64rW37fuv/9Ev33vyzLkfW1pZvZcdFrYaRym8LsIfKca5wRImQ0nhTeboqA+ML9S89qyXYhjOoQsaztzHgDGOujWpzvxQVzR0uQq9K54eBsRvCsygI54z0MA5+AQkgJZ19O4KUA72BZgE1Cyragr6CCCZ+ll1bF3pqdeCcC7rhAQ8qI/ZQG+aJ29hZNMb+HbXyj7OA2ws8cADX0hffvCB0Dt3cnRziHZnGN+tvnTJpZelyy67POs0YEfEGIvWpWdfmYOYzosAJF2AX5fb0esKTMn9t2m943ZsG07vfPut6cEvP5qOHT3Oitd2zJ0ABYI3SyoDOmoX4U/6AejZAR/HjxBEPLdPq/KhfKKM7bOcFA8lg5gbkH9h5kIaZ5nn7pFm6rDjaCyxpLxLAH0vDODtpPedgIa6WLx1HDdlGmOJTkS8Q9pzfMnE844Bki2VJoafG5/LZpXk35TfIxbKvEa+M9c+yTqPBM19+QUxMso4kx3lApjhUhomKQeoqoZKGnry5viaH88ExZB9uTYWmO9PD+ONuZvohamFdBJw7DxY1c6Lr06vv+c9aWTzLlwJ28gVYIxxb/KOM2Zb6GG0LkvEBoOLhcVemp2bQwfwToQ3PSSVq/yrSy08Ei8QpP/hh76Kp9lcAEzOqV5XQBWdoc7o6Fi6/Q1viPemsdME8My3p6Fj8KvXpKKP97CdVb8ZB4FC+bJc4c/r8DSM+v6gHjwpcj2NIylAUrRSXVswt0lDCNXyzkt1I2anc89MCnlpf/NocE3KPGRiAWxzKfDl8kkBUPmQrnnqRE7Q9x6ezXGXS+mWpB4GGEqebRrzz6f+zvB94HsOzan6ld8jMMKY8V6g3ZHRsdXNW7alTQT0dymrYOTg8AjLp0dwTmYLXQIzIu9NeP1t4p24CLGTXE/R7eH24ODYm+5+c+Oxxx6fn566IEhGy3HYcHW9zmvhuT7XEvh2S6Ca5d9uNur2awnUEqglUEuglkAtgVoC/78lEF/b2BBu4dg+ceZ896sPfmnqbfe+/ekFdtfCHBnBKJrg23wQUAB8AC8hXGEwNrBNNIx75Aoi8P1OIY1FbQ2fhXXF17+GiXl6npjCeOW5Zf3kL4aLZcwoHiRhGFnAbOkFDqNBbFvkQU+grJ8VK+ZGk/wIcMznFAtDVTBMA9b2aEQjL+pDp8XyMDuCtxCkADagB1A298zho0//0cc++RU6eyEKi/zAKofm2ndsCjnai2+UKpmvFzFjvdveQcKT6JAIB+5F7krYbL3mtjuu+uDP/sI9U7NLP7DS13cPtnfHQOIYhLOYlHomNhlvPcbARoAoYtCpGvpAK9xroJZkvrolywE8gV4IUmngBkpBfgYpGFeBLZ9VdQRCratHTfb08trnmb5t6w0kOOD1snHqSKHLtkM92y/eToJh1pc/z9mDBp0C1PBeqZiXdVE+BZT1GsPDimOw00rzs5Pp937/dwOEclmc4K6Ahl5Fw8Nj6dprr0sX7byIviBWgbYq5flFH6FpzKjwREK4gmTGUBMkcTdD5ZeXs8EXOs8Kr3TLzTek5w4dToeOHImA7QV0K+AOPYauDSlT+5Pn85qnHk/sn/M1j0WlQMjOKspTwEjZCza28CJr9ubSgc1DxCGjyEo3wJOWu84yv2zK8XNcgi73yt/rrAfIDh4El5QnhCnhKZ8FJ2xQGtYz13qlbrn2XOpabm3cGacoAw3zuQn6EK3oOW7KoaLpNWUihhglbdFq4SVLfvEQ854BiLrS9QhwDP1ys4Y5AK2z0/Pp+Pm5lDrj6TW33ZUuu/YmNlsYIfj+QOoqROi5xFfdsH1T8MgZLiIovztYdln4vsRulfIpMGMXBvAc1OtRDl2CqQeZQJmArzwuLRmk3zFkDiD7N971ppB58YCzrei3xEgFKF7Tgypf/Y7njJFJ2Tiq5b1rnnNEPYqSlboUeZY69iv0yVeLoqOweTFutlVdx7hxHf84Q1gSUS7Pi7gN/bDuxrxow1dUpStK0f6bKraq3lQ04Lnw4Nm0BphRI3izr7SjXEp7+XeRrEGbxviDTWNoeJil0hNp0/gEeQL+uI8NtHnv9beR8yi/kcaWFpeYurha4kxLa6tz83Ndfv/03vTmNzceeOD+5tzMnB3e6E2mYDKz9c9aAi8jCeRZ9TJiqGallkAtgVoCtQRqCdQSqCXwN5FAfNA/zyRYq6UzBR/iLLc8ez7dd99n59/zPd/DNntpEgN8M/V289fzFgY/Nrj7wWlJYAJhECxj/JWPdo1u29DQynkYT2E0aJqQo9Gh4cm1z/XW0PvGDEGsMLYrw8Q86cVDmjMFbZ+H0eMnmZTyX/zjSsOKPA3Bbm8RLrMxa7uCB1GfdjW8NegD7GgOkM1SSwEQLFM2IOsePXnm6Y989OP3w/NZCJoKWmE3vqPT3968WquhcKvkgICK9TeXAhxjId11b3zz9T/04z/zvXPzy9+PatwE6NOPF6IAFB6KmqgE3mEppQZsjAPAgV5BriaK5XsV5dKaZeLQ/KZl8QONZPVHLKIAYY635eKeMmiD40heqChGqQAZHh60pebZvocaqV64e+aqNigWuo6SKC/ggAAFRVDQJt1kdzpqogTkl/rlbMwv9Ta81OAjPGk4xxJidZx6m7eMA0aspI/+8R+mY8eOBT/h1cgzvX7s/8GDl6eLD14W8aHsq23Lg0BSJO6dV6p/F5nNA5TolSdIZj860AkvLeqq1y6LFEQZGeyku++8Np06M5mefvop+maM8LzEMOYRjTFLEC6HE5KzXjPBOGdlL8CiXHhKNhnMr+goOQF04zlmdeONDeJJtjo3lXYON9KWYeK5AZjpS4TkkSNzDoIBlgQICC2gAX46cDGOjlsZe8daOXsveQs6b/O9uELmJ8rLAEcAM5bnmXKRnjRi/kMvg32UDT7WAZFQKspn2VtZudrn3Lb1PQpNx0KgckX5q5D8z++9fF5awjORvs3Ozqfp2cV0/MIMXmONdNGl16Xrbr8nTVx0IC2zrHbZOWD3Ged4LyGj4A2C6nSeOQCG6KaHu/IKki7MAXjBg/0NsBV5Gg/OZZYLeI49+uhjtM3OiNBRF7sAZI6doF1ncCjd8cY72ZGR9uP9bSnGOMa/zJH8Hrd9ep1lDT/lHZ0BaeQk74pLXuS3HJHvcyWYx8kyWe8RVuTG45CpbZgQcZZx3OlRplOv80k6alE+Yi5uuHeOl7atWuYn7ESKeuiCrYROea549d5kfV/wUYaW/P1mffMzsOY5lw3gzrIVffsj787XosOM52q73SG24CY8y0bCW5Y/GOCU19e/1O21ebZtamp6D3rTofrZ/lb/MfRrYWW5N3jnXXcPP/HkE43J8xeIg7m2eLXiWA7rVEvg5SOBGiB7+YxFzUktgVoCtQRqCdQSqCXwTZAABoB/wPfQBWHw7IWp7ufv++zC97/3B57BEOktLiyM4AazGWNsBCtAVyBWAjX1JOMSs1FbTtMFAnrkaFCYNBQ0GjVs/JctqWxkaoZotBTDwuUr5bM/GyHVXWX42EjQjFpQI98Ka7Q17jgspRHmUktTgB6VWYH1sm7gYPxgLEPGJTOrK3hiEMscgKzd7n/imeee+uOPffI+jKXTQSTLJchV96/IE+OKdYiFiHXc12p3V5cZg0ar/wc/+LOvu+fe73vPfHf5e4FDrmeZVP/Sco9QV8uL1kEHWC8ooMoyMfSjJJfLmRfGtcOlFjFWAhEmn6lK6pPHRiPYcjnlM0NJGcAxxjUqUVcwxCVi0mnhaVO8lKJNwQ/aAe8NMsuG/SGpT8GP7Qk6GCyd+oIXHkFTuhze+6zwhbtUxlkEhbBpN42Ppk0ErH/yiUfT//47v5UefOD+0EeBF73GNP41tAU+9u7Zk0ZHRhQtoB6gXHg3yhHeVQBQJueSotFTyx0K1XY9yNqUbcojPGWaWQSrgDfMQPLb6ZpXX06dbvrKw4+wlBjXLjzfaAyqGvZ5vmRJ0oCADynPz7jMc4028jzkecwvQAvalMYKMf0EZ1rIbWV+Ko025tOeraNpkGaagC96uLmssY3XnN6c8uo4VdM05rOyVD/KOMlFHisBGugGCCM/+V5eHK+cw0/KlCRwZHl5K0laJRW6oQMKVVrW53/QRTeVS6nfZazkx6V5yidoc3ZHz4g3xhiqt46HfRDAnJlfSmcvzKbTxBpb6WxKB/EYu+Sa16V+dhldRvYuF/ftaGrqYQe4En2P/kVryCW/swRCPRYYw7m5eYL0C+DBXbwfsweZMhUsk//nnjuUTp486ZSKzQPUC/UmALLOYLrzrjcFEBxdpH2XX1rP92HIuRJVyKKSa8jHNrkv80/AU1k6DuaXw3qlbtSLXvIDfvK98rVMfhBQJPXX6oS087OgWdE3p7SR9SG3L92N4/u8Nq1T1XPOlDak9cIU3m9kwkqWLfz5Pih8lzakV8CxoiWhUxa1LgegWrDKuDZAwwDKxhqjo6P2bJU3aJMx6bAb6Tb0h10u+5Z4d83yngL/7DpFVogTt3rmzPn+40eO+HJaBUSF9fz7lNs11l/Y17UH9UUtgZdIAv4WqFMtgVoCtQRqCdQSqCVQS+C7RgLxFc/Xvt/1dCq+9wHJVj/0od/vvv1tb3uaXbZm5udmt+ApsZ/nTQ1BsCRCHS2vYOBjKzX6NAz9K38rloYJelBS64cjljdiqRm/KGK5cB1AiWc9BHS7waLQeBMwiE9/OQnwohjGZmSS8qvXhmXDUOORBlZl1eQz7Vomgy3GiAGjweTXAOzj2rY0hihsvB/NGgCyRj9UBr7wxQee/OSnP/+XZJ6MRjNAJlvr6E714Dv9FGL+xp3Igo8yWsIgHQND3aHRreld3/P+9A//8a/eum//wffOLS29A1+xq3U/6qEHOBuycSXWPcAYZ1Zgafw6NIIsEsvGcOwACFmXOzI8nDUABSuyhZ7BEpfgVRa7NRl/TfJsrFZeQY6l+Rn4DOzHOnqOWc5liFAPAMGzRrJpNTxTaN9eqjMcAaqqF+iydT3ag4BQ0oNOk3YEJgTG3DkQzw/ABu7d7RLdahJq6Oy5U+mzn/1P6X/77X+f/sOHfz+dPg1YoZ5Xbci/4JteP92lxfTQVx5MX3nwfjzMDgOAzMCMSyTZDZKlWjlOmgAGVjPgC0G9mUcstcRDrD2A8wmyynNiJbXZbEKgRMBQ0MX2ugRnZyu9dNstB9PiUl96/MknwTU7WtwBksT8LKPMnHFsQhwAKtbXI08giJvqoITjwS2iiOQcNn6Z8ciaK4upszyXLpoYSaNt5MXYNgXHkJ2x4eTNsYlxDvlCBELKfgBvvUI0SNuG/yhXxj3YiLHO7wrHIhh2XPJF8O37IdNAn6gfCe85miHFj6opxt0sO0P/BUTkxXLm+66Sjss+5cH4eBFrjHzHLoNivQiCvwRwOYPX2IXpmXRm2lhj/WnTrkvS1TfdkXYcuJxYcCMJP8pYWqunnh60ymIQ0Kp4gmVgTnZ8nr3fAiBzaaXeY3iuLRGLTN4CoKJc6KW6ic4qg8cefyKdOnWKPmRPN0AX9BNaTLM2u2S+4c474z3oO9K+utQylomGGOhtTAh7nYFDZkEII4PBGYwKb0Dajnnou5oxtkYpk6VnHxhbH3DObagrPI0OCOHaBs8jZT0wFhn/8/ubhxFbMuRFoaCV2xHEjnuzg4jLKKsCVV7k88xR9lp+c9nsCJlfNZkHecplZMb+5PmvjrlMMjMt4SyDoMWt7ymTbStPWfHseMS7i0b8XTU0OIxH6QTvk06DAP5piDnO76KR+bm5bTzexK+gFebbJK/OGX+13nLLrSMHL7+yfckll/aefvoZcNp4D0jdTtaplsDLQgI1QPayGIaaiVoCtQRqCdQSqCVQS+CbL4EIW43pws6CeJIBFHT/9ON/srRj587Du/buXV6Yn9e8aPIRz65cqYOxI6CktYH3WUMLWoMGO0xDjA/5ikENNo0NjTUNLY1Lje7iAaBBojGhseFn/wrGlqat5QtQUsqU+zBCpKoVJe2M6/ETc0sDV0sQutEGRrdeOmHEAApo3fAojK9+8B7SMn/lp7VVsIVm+upjTzz5qc984VPI4IQPSRayoe9KgMwOfuPEwAAxoBYgoJ1ua3A0/S+/9X+OXn3d6954fmr2e+eWeveCj161ghXZIyo1yyZxkCI43KqAo46JCK9SBsfRI6uNVLOxGlkW4rBoXtLkEAqOOWbqQs5XT9SPTAu2LO+9+WHtZvBTEAdPDWjBeQWcFeO4nDMv6kK22A2qrREf/EDXuE56f8iPgFN4PmEEy5M0mizhNP7T4HAnzbK07VN/8efpwx/+UPrDj/yH9IXPfy5NTp3HKG4TGH0UugBqACF6IWkcu/xKXRTAarYEe1jTzA6Ejz36aLr/i/cTzP9LASDrWTY2OpIEX9y9sgdYpReRxrj63XKTCmoL1ClZl17qOSceF+ARZUBvmBOtdO3VBygxkO7/8sM4kbEcUpHzD+nFnAmPMMuTpxDK8tcoQ3+LvNZcv5QbKXgBCCOaH9Q5E4dsx8Rw2oEHXeotpA7gDBGYkB80bRTays/5Fsm2zKO+74AyPvlhcBPPs3dfvi/P4ixQAt/2wyQt3xFryUvy+JGzaCQDUfl+rWzUyXI1z38CZHEN/R6HMvcd1nNXSg6fC5IZH2x2fjGdn55Lp2cWUrc1mg6+5ua094rXpMHx7anZwREXUBRPVd+i0UcBzVga6WAhS4YtgFix5ZAHZ0F+AaMl2pxngwY3aVgGLLNNuyQ4Zsw9wdm2ACNEjh09lo4cPRp9FGC1H+5kafcEyN7y1rcFXQFi+xZ/sAgRvUAezD+TuZZznOVLcMzkOOWU3980E8kg/w7kGnhblbJupKqcYGMZK8/ld4JtmXKbzuuqHnmW23iUMjmv1Mkme6FTaHm2XDkrb3m2tagPz3o6+s8U+igv1rHdqpz9lnbhIwrzw7ycX8nGuio0/32HSBfQrDHI0uex8fEewOgyQHhrbn5+YrnX27G02MXJEiieXS+R3SCezY1du3Yv3XzzrUuddrv7xc/dRyv+0sv8lXbrcy2Bb6cEaoDs2yn9uu1aArUEagnUEqglUEvg7ygBDRk/7/+6D+tsBFhQ05e/mq9+/C8+s/Sxj/3Jc9u37Xh225btF4gl1Fnqrm4lVtOAxgAG2LIeZRhyru9paMTqJSIFHInIwqjUEJIDiXoBHxonGvKW08A329vKJqMej/ihMbJuOGGcRl1LW9V7dmGrDFcrheGroV1RlUbUx4jWYBPcEAoUUAkcjQBROkbxrL8zOJhOnD77yB/92X/6JEW+6z3IQogv/iMLGOiJxPdvH5b9QHfvJa9O//o3/9cxduR75/nJ6R/BTn/TwmJ3f3d5tU8QEs+WZW1MvCKMueNoOiRVXCsMYEYlDE0zSY4LPymTjU3aibER8IqdC6Hg+GfPMOP7ZLb8KfhFUzGO0gqPQOjpVWI5VVBDPrypABEoHl5c2bMqq6HgQ66bP/EFlzJPUMagXQOb0BkD9aufRR/Z9TRAhmcOPZv+4CMfJgD//0Xsp4doG4Co3WInu/G046Ldaf/+S9KVV11DEP7XpGuueU264YYb05YtW8PMHWKHuxZeYHo1NvVGA+AQlHNeXDh/Dq+yB9IXMIpPnToRYFynMxS7GM7gnaR09YiMDQnsnLKm/wImIXRkrYebYHUADM6zXiNdd+0+6g6kRx95DLDN+cK48Izq2fYWbOLa+RFj5w+fmdx4oFx77xhwn0fasYQnyiwvTKeRTl/ahRcZ2xAA3OgdBl3aCS87x1SeqexYRdw3znk0zIYoMrA/keIdUeWTEXOXIg031pWMLFJHCEL27K9nOyDNoMeFXqzcpbxk0jL53WDReEdU53ir0Hb2FMs7UepZ2MNrT5oLLnNcWooYZD28umZnZ4g1tpBOXZhO071mGtt9SbrqpjemPQevSa2RzQCoY4zvAAqZPYrctCAC6yMTdaqAcNEDWOQthe5mDz/bXSRWmDtYLtJmAcjkV69GPZQ8BHIHBN/Q1cOHD6XDRw/H8kr51INMLz/BMnXvDW94I/3III90PNbek8hOfkJmytOxgCfPiDpkW3aBDDCJsWEUQt6WyfXy2fdtJGlsSMo3j0zOtFwGphkR9a1KBYgyJ3KlUx32M8aZe8uZnLOO7wuTQLvgnqSl77shbqqCcm/WGpuUC9ootiCz4LXjVFjLfcyVvZZm4cFcRJv1Eqq+Y5zPPg95UN65TmzDVeZ/A+CrT88yllC28cIeZ43lPuRzAB3vwMY5YsadIVbZ8oXJC32f/8xnlsl3sGwlM1D/rCXwbZZA/u35bWaibr6WQC2BWgK1BGoJ1BKoJfC3k0AxGsIy+LpVNWswibR3tUwbhOV3h8ve/GJv8bOfv//Q6ePHz956662z/a3WFMt+tK4HMQ6GMLADvQCcciUKSy/D4AxzNBoDGdNzxMNv+zAwMBTCKK2skmIYeS4GSDE+zCvPI48/oltXNvNZ4yV7ekguHmn0YHjZXhh0Gtnca6gIpgikSIF7rRvZBDtrLs8sLT30Rx/7k79Y6q0WgEw3F62R7zoPMjv9DZJmHtLUUbDV3XfF1emf/vNf3zI1u/C2qZm59yOttyx0l7ezS18fw7HcXUI8IDaMB7Yl/1UlCMR4IuuN46pBbVo1/jRN5DvuUam4I8Nx1qj37JhlA7PBMt78OR4AS5SOwkE/8iBp3C6L5aVn2bsmgFFoyUcTIEp6tu05e+Ooj1mvwrOFfHaZo5sutaQc9AI0gu8BPH8OHXou/e7v/W76xCc+nk6ePZ42jenpNRTAx6ZN48Qf25S2bd0WQdENhj7FsrtZgK1z58+m6ZnpMLznCbauTtpOpz2Ed8+ASsiSRCSEvg5jOC92F9ORw0fS/fd/MZ05ey4NDg3BiHGnDMzfoo/G93L5J7xmj0jObqABmEM5Y4PFHGFSuNSRxZ3p8iv2MAda6cGvfIV6eJJRDmEHKBCVvHcSA844gey3fOmZ6bVyi8Nnlq3mVpSlDKtMU1qaT/u2j6URZo9eZR3ODZ4FqFMAA2lZncNx5me0Y9vBc9BXBzIIFO8Anlk2eI63lLWpqSpBKWtdvH+yzvCsAKE2xBsDQId4Z/As31FXerQlIGe7XAVIZH+8d0l2nAHD9BoTdHLJpR6HenWdn1lMF/Dw67XH0oGrb0iX3XBbGt22O3apBHVHz9H/qm/qpPrkXwsct6LfeX74PsrLLmk62ojNGGjHwP9z7FDZXRKoY0k7PEknA6QVUEo76sGJUyfTk08+CTgKv/Dp0nZ6Enq+ddv29Prb7wivNPU++m3fOeSlHEE/kCQkVD0LtpUVWepDuY/Yf+RZ11TOjoh0OK2laK+6s5z3Xy9tfO48tWx5D1hHEOsbpZjjUaD0TXnTHv/XeczX5d5zuVY9BcgcJ3XCjpRnpd3Shv2MOQKP/osxpuvBL/eFbq4fMuRXUF/fQLuzOjIyvDrOOwMP3FH6tBP9ehWAPFO8xbanaQFArW/njh3EtDs/f+TZZ1z7TLYwXJ1qCXz7JZB/I3/7+ag5qCVQS6CWQC2BWgK1BGoJrElAwMF/fja/eKoMCQ0KPvb90M/Heg0/3POnfX7kH8816igZhTSGDh87MfPnf/7nT91yyy0Pbtuy5RTBzUcwIPZgfjXdOY8ljysYkCsY9Rn6kCaJnwGUCIDohmDssTC6aEojR+MtdsuzDxpMABVyKD/BF4aepcKeXWc5ABW5NCA5BMI41uSNFqkBmWiPnyQMHQ9lQGegi93az/rQMLxYHugGnQOT+/Zf8qWf/c9//jOHDh8+9ehjT1gRR6Qwu7M1bc4rIgkJGdRooHfZa29N/+Jf/+bmw0dPfv98t/ujjebATYBj4z2AH8FHdlYUfWSMPZA/YIuWpWMWScOWO4FJQQjFqQHpdeiuxSgjeKFBGmOlsR9Hjl1ltuCKWhGx5LwOwzWPdyzXc5hox3p6bag7tiMoEcCT4AMH2TQnEGJbpuzBYn/02Am94Zn6ZzMhiYpel4D0H//Ef0wf/Y9/hOcQnlKjg7EEcmW1B3/9yIKld4BTs8QKewqQ4sknHk/P4WV24uTxdPbMmTTFMsrTp0+ns2fP4iV2IZZN9rEb5iLxrGbn5gLwcAlyG2/GLvwY2y/vUNgCYJtMJ44fC9N4YvOEu+NlA5xuLOO55dSW5/AaA3QT0ArvMGTrvJKOyy07nG+5cTfSHkoPP/Iw8JW+V8rWAxkq7GpMlI5jE6mat/FmsAzjpwgbAJKcbJkfBuUHlOuyzHKkkzYPtVInEQdN+ckj5eTTd4DgXiQzeOKIODh6UsVsjfEVSKqAlmoMrONQr4htU9K+BV1RM/57L2C+QiH/RdnIg0PPwWeobABhqyx/9d3iO0igg+VuoZt5LAGjeCiYVMCxRQAqgbGZhYV0ll0qp3p9qbN1X3o6yoQjAAAgAElEQVTtHW9Ley67NrXHtoJMskMpR25P0Nb4YCbahyG1S6Cuj9XI5gXgRBl1HBYzL3EGHOP9hqcmOkIMMpZxFoDMnUuNr0ex1GFXSudOC89Gd0t98qmnCOq/QP8E08T26QMunzsv2pluuvnW0HPrxbvSuVDJh6zou7zGXIXTAGy5d2QKWOlz/5QSnpte+8bneQGMnHtRg7NPIvmbgBvH2aFae6AuWb4qaF0PecqgE2qLDLw2v5yjhapc1ULU8Tq37yt7rfV4FwRt30NwkXXMtuXId48VKe9Bjv9KXh4vJeBz/m84rOb7xvdGjKOMcV1kIejpiFs3dJX24/eQSmdd5kGz3UybJyb6Yul1YG39w6SR9tDQEM7NiLkxe8MNr5v+4pe+ND89ed5qtCKfL55y/1/8WZ1bS+CbKYEaIPtmSrOmVUuglkAtgVoCtQRqCXxTJFB9en9dWho1L/7B/OIf2Hz8xyc+T/mC57MeGwlbZYBMNtBbnP2LT33q1NFjJw6Pb9ncHR0bXV5cnNfoa/et9g9h0vcDhLHEjnU6ORHEnxhIGDjxV3WMAndN4yd2CJ4aWBURLJqP/Wwwri/x0bgMW6UyBPTwMWnEhqERJocggkuCqvwwG+iAGSRIxDPLh1Finv+4J2QaNhKhsrE/lpZXu53B0aPN9vADu3bv/dLIpk2n/+/f+5AkKBFcZGvGnO/CVInLnmXBAVIQqGp5y65XpV//jd8afPbI8bcQXOzHgCvuZp+14aWu/jMNHJVW/D7GRjQYPzLG+HOYvGZg4+xYeLh0KxuNWf7FgCzBwh3dTKMYwtlzKe/yl0EUDdA1FmE105DlPDw0j5Fqe3DE8IZnFXXijKFqeQ/pyKKsZ33K3Y7lbqFvGUDRqBW0aGPAPvPs0+mPP/qH6VnOLpPr4PE1SEwn21siPtj58+fTzMxMgGCn8OJZAkTZmBqAIe5w6E6VgwBgW7ZsS7t270vj4xN4g3XSPJ5JFyYnocESSiadu28KfOTlfC7vYxkrZYaJSzY7N5t2bN8RgFqZ30Xn6VAMojtchlyq8cj9dbkjY9Frpcsv3w3w0Je+/NAjscwzxsyxirFjTgGyRVKYJmWq3JwOlIn2Ig8ZAsS4RFT5CzwQtDBtwX1s28hA2tymL6tLLCsDN4rxC8EHQCYNwYMYj9xK1DffwznvOOZyWW/s7zqvVpKf+B/vC0pFXm4lP7YHcQ/fax5l5MV4ozqelW/2qvJdoodYBsyWAvTMSxwXDJQPWDbLksdTk/NpZrmZ9l15fbrihtvxGtuTVlrDiZD4eKhVMqMN9S36w7VcBAhGmxkkUYervgJVCjoJ1sRYwbAuuYu0uQhANh9x6IhBxrtUeoJj1m3hsmcbAqDK8TRA7FMAZOxADB11ZjHOynLvvlelW269NWLfGRcv6/76PI179Qf68upZPgWKlHtsSPGC/gggm/ISR8uVvtMXO8KtZ9vXly2uuYdqBsqoG+Uo6nm9fpXPc/tlX+2nyTJr4Jz8VUd5Jh3Ll7RO0/dEbkM9NV8Zlecbz7ZZUuQzNnGmzvNSKJZzA1Cadgv9Mu7K1FT4Cd7kN/LslL+DmjiqNVaIV7g8MrqpMTo8PMSvp614l22CD3Hged5h87yHFh74/H28WGyoajgkHE2s/Sj9WMuoL2oJfIskUP2W+BZRr8nWEqglUEuglkAtgVoCtQT+jhLIn9v5g3nts7milT/as1Hhs1gqFt/X2dgo4EL57MeOWSPBZXzKa0O6IMdVV1PE4vnDT3zy1Ec+8cmP/OB77n3kAz/8/hu78zNvYxnQndAaAjcxbL/L7voH8C5pckhQDwyBhQigTuz78OLhr/d+zGOiwRjXGEAaJrGzITyGacE5GzwaxuseJXKm8RH1K+NL2z0b0Bo+leHk2b/i22dSeNVgXehtgcFGFWyUZotetc4PNjvTM3NdbFis+rB0KPIKSJVolCVCDnks79h7RfpXv/Hvxo6dPHU3hvp7G/2t6xJRcBbmjYHVxwrJDGz0EOsKPwxiXoy2PC56SpADIOq4GDcsj4A6yJXtIPsVxjEMXwCJMkbqQATZ57l1XeZk8CCfm+8Y5oER8PKqAF3F2M9AmMZ71g/yHWm1WZ74IaAjv9bHeSdANGOAOR/wigvdcnnd5ORceujhZ9IXvvA59iloEXR/JPggfpBKnowJJnBF/CDqQpFJMgKINTQ0Apg1ynLLibR58+a0edO2NDExkbZu3gLw1aHMaIAwgjKzs7Pp+IlT6eSp4+mRR75KoPXD6fyFqTQ6NkwMq2HiXs0F+Gb/WWYVPlZHjxxKBy+9HA8U5ILo9XiK9pkLKu8i826QtY3Gc1sCpJ5m0wADxI8ssAPmMJ5kY5vST7/v9vTEM8+mz3zlKRwoxwOQiTESzXKyS0iBxUwUXHKOMpfiX8xOZMFzvAZjzPo68KEn3FA6en4hXdjGMtE2Y6PcBV1JfTom0kiAMfRHIM75HzG/IMV2GdGsa3fVizJuAqne6xClmjYYm+A1eDGvETqYtQxClDcFLCOPJnWQPpS2cyZgmN5trFoLwAwAyrNgjmfAYILks3Mo8p1nKfH0IscSMd624DV2421p1/4r0iq6tAjg5FxwIwV5cU5lfaNvvqcCZMrvLIHC0HXeeeU9hQSDHfOtS+3oA9tesLSSty9nyywThiq8wphcmb66nN/l0S+k6R8hlBt/qoj+s+lw6PxwbBhR+q8sbEvZlPmTaUonOHDOxBxy3lHO8a/65TL14JEW5MP3d6QNq/9CDjy3HcRD9XxtB5dL+VwryngpO5bXI85z7pn1cr4eotFeVS///cJn+XeB4xYKlH9QVmFCBx5Db+Q1NC6XL3KvyK3RVgYh36rdtfGDwdx+lt9av1FMea2kEDHqpOm7LuhE+6UuEkdnchvyh2NofwtOWVo9OrI6ODzU2LS8ebjXXdqPp+pCf2Nglhh4CxfvP+Cyyzna7DqfkA+dUbJ2ej0ptzrVEngpJFADZC+FlOs2agnUEqglUEuglkAtgb+VBDAdMAX8Rv7GKUAni+DJUgyMv8GHNEU0zda+wNtzuJ1wP0/W2d/9gz8+e/jZ54786q/8d5Mz5yfPrfQWbsUQ2YcxMWAAa201/G/gcJn9u6Dh57yGrcY3qMRqo4snAEHyXSqEMdo30IcxuBCGvAarZTWXNW40Vk1hNGMA+CxwFq6jPzClvQA0EkZqGNMYZHoaRJtVOYEdkRvosRqw2cDWhTvi0DcHG2B6IwPtwZ3Dw6PGIDsLYSzTNeEqZEXxXZuQH6rU34+Nv/xzv/CL6dz0whXd1fQuBHUPw7ll0SBImMiIXlgm5B2gCQPuGCjnjck8bbWiZxHDCnEqRMGx0N0ok8UqeOq4mazrdTli2MI4rgzkim5WC3Qhqq3X1TDdOO6hI9CVQ5dDYk/Hcz1vbEOgSq+wbtddIvP9CksqH33s4fTMM08QT8zdJwHQMGP9N0kg/aWFuVjKpom6besOgvNvlnUAInbAJAD/9p0XpcsuvSJt3bo1jY2MhxzkQ0DNJW9Og5gKrcF00UV707YdO9O+V10CUHY0PfnoY+npJx9PcwSA1xusMQhQglfa2dOnIii7gNTOnTu5JtA//NpXQRxjkwnsWa/ZN8g0y/GR7CfjFx5uHQE9jvHWtvQLP/H30uS//M301WdPETBslIEh9KAOawBh/SzjY2/S6BMTKc+zfOegKkhOAAl4u+FUGO22mEtLjVY6R8ysC4u8KPA1XGanzh7AuQsNW/DqXA5d4TroQDPGyqnJddYXp1vO92wfzQ8MV3g0qwxPvMhTUzjIa3mybNE7y0jXpZ22Y7nyvPDiUkurC+Sb2JAVPgF+0YtFjnlUf2ZxlT8QNNLOfZemK298QxrZvJMFpAIdjbQAxK6OCuTCZMgqdE45ce/UaDJrfJz7IZ/53VX4tHw+LAO/yjQr+JrMnle2mi8bvWsDqAwALteVnl5zfepk7Mqa50ihE/KAuXJP8eBBGQT/a2fnWNaBkl/KlLrem6SJX9TadVxUP+wXlNfa887y0g5QM55nGfmsjLvn0r7tRXmeO9amNR4cg433XGeZZtnaTAYF830UrsqXfhX6ntfyqoLlHirWglYlJy4ybF/JqAL4LOPvrxemNX55AE09mZlzbgSdx6eHnuE1NsL4H1jpLk03O/2nr3r1NUf3H7z03LNPPnZ2Q/1KYi9sob6vJfCtl0Ce5d/6duoWagnUEqglUEuglkAtgVoCXyMBP7G/9jN7PY/P/fj3wq9lDUpTPkPBL3oPoQIfvbCChV88BQsU1zeD/5mboydPz3/izz5x6J33vv1hDPlplmHuAozb7gc8BmnXP+CvdLt9xszpEXRcoC4Cfms4AIIF/hQ8YaRhwBZPIz1EsDEwngTGJAK/Gr7cC63EdRjCekT413sMjCivQaIxbTxjyga3GMYYvII5LgXSOwFbhFVvrcY8qwRbg+OrndHx3sDg4CLhkeexZyZ/49/+m/M0xF/qo5/+8KDh78xUOvC13KsE5SnuKY3W8qbd+1rvee/7XnVuauYeHGjegfG/3xhdAAFLyA/7sq9fsQo0aNDpsZKXEJHpgHM4jiZtQwElwTHLBqDCQBVD0zELocoCqRU7/rlkjCV7AQA4XnmJlXXUl6AXY6wBG7XhLe+SWGxRg/VnsAAvRrw1ApzjocstDeRlOflxSaEUXT62gieR4JWxwpZYOnz08LPp6JFn0Z2lWBopYKY31xxLKRc5qxub8Ai75prr0q6L9sTyxxF2LdzK8smrr351uu41r0379u0jCD+gEx2V9hzLD405tsSSuQx+VGAcAl0ChQSTiRhk+/bsTbt27U5Tk1O4b66kCQJ5Ly6ybI5+yoPL8VzWtXvvXgBlZAsgoQyURpYIAAv6LlinLLOXkXMDLyTmyxLLPY1ztn3LSLr5phvTX3760+zGOM+SvRGeO1bF9IEashLwiCGKa+gwn2M8kF/sKqiHH+23WS7a57wE6B7vACYNrqRNrPZ0SWADryHHBOJwGdTIYwzk2XFgXgpfOXYRs5D8XBLwwecMmroWuoO8/CcdvYYEqWIkKcNsD3rW8fCfsvY94VkQzKWKHvLcBQBbAuAiUHrs+qhsjP0liOmYzOHBdX6e+p2xdBXLKS8nLl9ndEvqMgYLIJwG0WfiwFcGX5+n+7625IyH+bk65zjl/gvM5bh6GRD2Xh4X4MHdK+fxWJs3QD8Tsdtbgt9MqzWQd8VsE+tMecUyYmR75mxeYunumjmOWjeeOYdec/316ZKDB1muuYAsfKXygxTvatr07DvX4RHIDK+reFcy/xwnDnVNqXsfYwmJeGb/+RfjaEerayRPnuAkUkBenOKI5aTcOy/sv2WyLpgXTGWKkiLpwVaApgIi5Se5rVwp45PqDJxG/cw3S1ud945SjIN1ohH+HqDeoHN4Nmbec36uH+zJ2Fo9x9K61goasst4+s4TlLe9WA4a8uIh+XIS7yCvkKc82Id4//jesb6yoJzxzJArvrrKHIy61ezgcbjI789TAPQn737LPTNPPfNc99jhw6LEaEv+F7xAoU61BF5KCZTfEi9lm3VbtQRqCdQSqCVQS6CWQC2BkICfzy+W8mf1+lM/25+f1p+ZX+74Rs83X1vh+dWff6dF5WHi26jR4bw8Mzc/e99nP33i3e9+10kCoQ9iyG3HIJ/AyG3hGaa9sErAqlXikTWaGkMYldkYwZQJ4yIbDMEblpKghc81XrXTNYq16ATHNAQKaBaeIlWPwkihLxpwPo+lfRqTuplVSc8hMjBQsEqwVBZZhzS73NcYmtjGlmLDA6tETMbA6Y2NjZ257/OfPXbouUNzmh8kvwO9WCdm7ndQil68KL/20IBTuPL1NZdZR5g++PO/uKPVGX3HSqP/+xa7y9cgTl2nkCvIEtY4Y4ONt9EYzoQ35mlABhhWGZel6dC7SoqWz+J1eLMXSQNDVsPbZWiePSwXxrnGpUZmdZ9pZl3R2FRnSoD+2IGSYdYwto50wiBlKAvNAI3UGUbXgOYCCnPzM2meJY/HjjyXjhw5RCynGXsOmMIOhoBmC/NzaX5OL7NmuuTiy9Itt92e9l98ELHoicaSRgC+3bv34Dl2WSLQdoAdiyxrXCROmYHTBWHkcyUAR+Je0W/jXGlYh4cThrJelRrom8bG05aJ8XSOHSwX5ucBuliOKHADry7j7MLTpVdeDqg1ENPIfgmuxNxBOPYpgELkJkCtoe7SO2ewQ7AE4NZgbm0aGU57X/WqdN/nPsdyQuciXp/OP8pot+PeAn3vyeFeucUzylA45qkUlbn0UZDUj9L0LU2ng9vZ4bMNAAFQ0nYMrAsN+2GKMQmlgAKyENAL+IhCjguMRDnbDn3hLnQFGuaBEESfHWN5FhTUo0rQQ086Hkd5r3srAkzVfSUnYyTq7Wozjr+gmWNCVprn+sIcseEAx0Z27EuXX39r2rbnkrQ6MJzYliEtgmayo2+AHvY9dpUM4EN9teUsK/voodycFzJle/IrEOmZ4a9SBsgMTK93IbsIw5fegQbcr/pGeQGyNjuq5t1W1+mfPXc2PfbYI7FsN8aQDgtMuaPlTTfdDOi6K7ziBP+kp4ecZ5PvzADF4E81UZ+CZ/qifiI5+KyAnSgvIJT7aX37bJsmT46znVWePssgWX5ugeh3Vf/5dR1r60oz60i8u7kv+lLqWk9gu8hYnTfPxj3HAesC6aVuPA/a8Bu/I/J7xfbk13dNDJN0KhrxpNDbkOdzk7qaeeLGttFHUwDwUd73lnqZ+ZAXk3pqvQBJzWO8lHvOkxXeKq3+HuEJzgw0WyfHNm06hyfpzF996pP4Z4bfY9CRUp1qCbzUEsha/FK3WrdXS6CWQC2BWgK1BGoJ1BJAAn7+fr1PYD/4/fB+8aTxkw0gn/tB7r0f4PGnfDMj+anzN/7c0X6SCmYm9inXzx07nd73Ix946uyFyd/ttEf+n75G63gf4ITGGW11McKWrWTcJoP2h6GPcaZRjFWKpxeGPcaq5433yxqvWooeGEKrePGs6EnBWYOuh3ePuwhGf+QIGnqwxO5rgGPmK5/wTLPPVVomj+WDq0Nj46v9naG+pdQ3Ssz5PSt9A5c3OyP7P/YnHx/54E9+sBTXCsqWUMn5Djvb8/XeP5958hESaNJqK91573vSRXsOXInJ9g68xu7CBBsCDmOZbV8Pww0Fwb0odCgb0HrotbAO2RI0DvFIZf/1UhiskNlorJrnfRzUz5imBqWgVgbMNBrzrn/SzmBIqRc0rVcNkXRMYT6Gt1jo4PPMyRhM9MEYXpZvoastwVV0cmFxlt0nn0qTF86G/sQyO8CxriAX3lstvHZuu/UN6U1330Ow+6sBsrbgYTaUBtpDLHvclfbvvxhaxChDajPTAGrUc3kjMoy27EubeGaePVz+GB5OGTMKfWU8sLP70r4DF6frr39tlBNIGyBwv3H9ZudmANzmwtttYJDNAgDABIfcVFRaJo30OXY+NLi8O3S6xC6GEAH3KCvYYX+mzp9OV+7bmX743W9NfQsXCCMIKOh8dG4io9gplrkWNBmr8OGs5pKyp1PxTOCuhz4wr1KX3TnPzC6lUzMLLEMcYAmioFM+5EWZW1cQVVAjwG6uA/yWf+Nn0cYK7w+nvkuuPcyzfwawDyCMc5SD1wAHLQyv8Rqh3CLvA4+ow3gECIYce3jxdQEIBZ4cXzda0MPPY8E4Y8jt9NRSml4dTLuufF265ta3pE0XXZx6zUH6359m5y3HW8N+4B3XT7B89/0wyY8JuB15A9JGtv3Ri81zVc7+Q82+KgufdXuLcS46LN/yJ8hUgv/7TF33fWpbpaxnAUZ1KssEGA/g1rwm46HXlu9T4llFGwUcC/q+i6EVcwleog3PtGMcO+d8PHOe0bA9iED50Qf4oA9waLdz2/RMnj0cJ3XTvsbBe1zPPghG+VInn92xMufbHoUolsddnmLczbXdkHPWJesKlOUa3uUkT3k0Ml/KzD71E2rAd4t0siz5nUE/i1ytHf3leTlXJNdOWUaC8tCm64x21lPrMseUEz/Eyzijp5yjPcrTFa7z2BXvNmVsnEBTeTfk8s1hxm9Xq93Z2d/o7zCerntG0UkMav6dHnf1j1oCL6kE8pv/JW2ybqyWQC2BWgK1BGoJ1BKoJfCNJcDne2UorJfzo/pbnLQ5tIYM4aVt0CFyz8gkgXp++Vd+7Svzvd4n+NJ/Jgw2vBxIK1yDphkQ3aUuVOZa+8Gzhri7UZaz17E7JTaAxnmAYQGOcY8BbL0wNK2DcR2GUUZVcj6G06rGEuU0eMLo0RDSKiFBgd3oMJYxXdvDY41VjEcYpEON8e5yY/9Sd+Ug6y93/vRP/2yUr35A7bspKQstX4PA9SPY5sJNd72l9e73vPcmFiS9Z6m3eqvL/bJBvwqemHWqGNFhHCIzzzlP41ovomzgZUlVRvXXMTI30rR8uZem19LynIGynKf+lOf5WR7XUlY68pON53INbYzXkuyT5UsfBJxokgNaFHvmqccIij9JJZa4sSmBSSh4fm4R4Gsw3XTjLemWm2/HG2cfwEObeF4a/800OjIRccdcJuqSPXekDE8g9Zk2BUICrKAxvY06g3gA0bb9kIJlBBy9L/GiBPl27d6d9u3fD38sUwb56QyxWyIgzyzebEePHg1AUsDN/khPMEJPNYGhBQLLz7B0coGdEAXp3CDA5Y7RZ8ZLoJqtaFN3+kK6+7Yb01tuvwG3JVYX9+YADDDgoYUwkV8e/5Aj9/LCgyxn7gVi6ECWFYBGk00KuniinWCTg7lVygIeGsGOmtE/+xH9jfEFuIFf+d84dj73EFAKDzDK+Nxy5heAJ8aHfgigC5bHOyVeT75fwBJ4Z0RZ+woNrz1LIwCzKtaYMccW8KCbItbYmRnAipFtxBp7Y9p7+WtTtznMusNhAvIztrw7mixbFdh0nBzT0EXGzuS1PArKx9gy7r51ik5axpzSV8/P6wv3JmUUfeE+yyGfg3bRX/Q1t5d/D6iv0hKMM1lPGk3ixLl7ai6LJ2LINdNbL5fHk1kX4FfxHpM/68VRvWe9Lvx7bVorU5WNTPXmBcBhKe/zwsdGWl6bLGdfC13zvTeVs9c+L/3N1/ArnwKPPBfIK7RKec9oW+R7bSo0vLb8C1PQkGI1Rzfy6VgLsFkmDpoXECvvJcuaL/hX+hRn2fSo2rMch43jnGd5wNdmc6h/oL2LPxDs5f03gWcqEyq3s4HHr2V4w8P6spbAt0ICeTZ+KyjXNGsJ1BKoJVBLoJZALYFaAn9HCYRhraFKfa9N5cPda7+a85dzNtLMe/H01z1/8Vrm+n3vn7Q9nj55Nv33/8M/OcEn/nN8zC+6cyW7//FBv9LvsqAVUReSRqUGiQBXeJXp+aGBiVFYQK8lvTyIZbTs0qcAwjBq7aWGfRjYQFoYERr59lnjmMoBjtlGPBNYC2MxG6jKqEvZucWVNDS6udHHjnv8WOYv9Csa+d2V1Z14ahxc6vYd6PZWN1feHgJEmXGRgsoUkf53ZsJg1NshfFuwnFNr9aqbbkvv/7GfuHh2offDiPp9qyv9WxCxUrTfbu9IyLjcX/stkBM2qNccBXAK45EattAEe9NwjNY8bzB2Vwja7hHjhrFu8roYmgJhG/VYj4/w+oBui+VsazS5l8ONnji2U7RZj5NQrQoQgKiWJ0f2TLNstBv8JuKOPZOOHz8Snom9FQO2E/AeL6v5OT0W+9Mb73hzuuct70h79giOtVgeqafMKsspR9P27dvT4MBgxK4STGMnV6hmo1kwZYSljG30fnCoTbyyQbzIBMlazAU9fjKgMc9SyuXKw6eAZO32YLrsiivTGPHOFgA/5gG6wHHC2+no4UMAXN00PDiURoYHwyPOtgRXegI/HHMs8ZzFI8rlgPZnmHLDADt6+g0gSxehOp4ri3Pph959b7rl2ktTo3uBBqaIH7gEwOTMJiG7mGNc6n2G6xR5nDlcstdg/rgrJTueBoi0BOXDZ6bxJGOZoICafDFWlV6FPhSAJMaMMQrdYnwKMKTGCYA7D0tZxysDW/THwfWIdwlvBz2kAPyIexhnZenyVmO+WUfwyA0F9GwysL7xw8x3t8pZPMf0Gju71J+2XXZduub1b0vjuy9NPd4RQ6NssoC80JwAxjoD7QCc1FOiGcZcsA8u8XU5oB6JpqzDmpHoGfWB3WjbWQVgojx54lGSgKj9VKf0QCxzwHORic9t13doxH9zLEj2U1313FXIuDb19K6Fp6Gh7N2oF98Cz13uq7ecPXL+OLdi7tKuY1DmhRtn4MwYqYxN3DD5zQ9PKZ+jAzYpbybr57PgVX73lr4UcFSZmMxfOxhw39GlrQCt4d8liMreXSytZfngkWf2MeSrjpBP5ThkIYBg6BXvLuWWecs8Rf9p0fak6Wu+tC1vJa15l9lnD8pJ37Im8/Sik/voOnxlmgK/mQ8d47IGKXOuOLw35bbzWHDLBfzhggYNOqRK9W+G911Q2MHBbhqJYJAhN5+vJ8llkut59VUtgW+RBJyLdaolUEuglkAtgVoCtQRqCdQS+FoJ4HNByB7yNREefebw4oNf+eohdoR8tq850CU+U5NrADKClff3rWqkmDRMTRpVSwBhXYL4a7SF8Yv3i15kXUAyg2oXD4tYtlIZNIIy1tUQKWfpFaNFbjSoDPBscpPGLkbJ2SkCpRuIvD2Kgekum03s0j7sUflY6p9fWNqDjX/Z1u279mKMdDA4NELsmldr5ocGyndSWpeLNmajab9BLeYuufq69HP/xX910cx87x2EGSP2WN8OjViWn81Rp8dh3DGPbJQjU43MYgRLNwzLShze+8xzkVGcMb495/JZjBuvC8hmnqmcNSKtVzw0yjNBpTDINSYrup5DFypeNNrNM8lTKVf0hSzAPfrSj9fQmVPp0UceClBWUEYAwnLqpHb/wf0wWZsAACAASURBVEsuT9de9zqWznVY4jhPvK7snaOH2+joaLWEkV0k0VvzBKpsU6DLQPmCOG1A4g7XTQzoAI/x+NIYtqxgQ9Fp25ROSSMAcFsI/j/IOdzceGCZyXPnWTLnjpUZuBkdHmGpZwZP9ENxc4UAfwDsJqfnWe7JDpqARPbNuGTKOGSBoPqYc63VxfTTP/r30lWvuogYYlMsjiSOmUoPSBamugAK4iwyDcHAi96fxk5zrjpR+vCig1qa7DbTyTkAn/5BPMgEMMCzmGe2a/+yt1MeM/ko41fOazHb6AvVg9cCFJUywVegoILrHrQnyChwzrXPpe1he9Z3aaVgkdXmADkvLCynk5MshW2NpoPX3ZIuu+7W1Dc8nlaanTS8aQsOsXnpou8uxygOATN4si+Os8Btm3ICj7alR5ptRb8oZ4pr9DGW/3JvH6zvYfLsDqLuoinI5XPfh9Yzec7Lc3Ob8mGZcp5hA4mlCtA038Ok95h6uJGO+UWWngt4FDwwRvaJFi0W9AuP3hfa5hWa5kdduiI9Uxlry5f6BTQubRceowI/LGfb9snrOJwmHKWsZ+doDGBVsdTL5XO/fXcUWnbHZybznG+M0BrN8sw+B43SNueN7fqs3EtrY1nvTRloyzzEcy49R7ucbcP3V6lrfqGpPM3nXgJRk8tRSm9rDXS2MzRj5AtLliTB3LGSU59rCbwEEshfci9BQ3UTtQRqCdQSqCVQS6CWQC2Bb5YE8if6+tdzuV/7nF7L+Ju36Me7qXzQl5qS0pzCbFk4dfbcCZYvnlhZnNm1iqUcy84W58FeME4IkI9ZEqCAHh/S8y//zTaARDEolzU+s2eShpvGhPHG9FrRsOoDwdJ80IgyuUslGA5XGbjJxgceB9VzC/fYsfL0+dl0HmP44qtelQbHJgi0jdFCQxolGinG+ZlbWByfnu0dHGi3DyCnQxBdEPDAE4IG6OHfQWby+K1MX886WmdVA0wOLMl6V+BB3B5m915+bfrFX/rlzbMLi98PFPI+PHVepXFuWeTeAihjg0eXIzIWDB4VAUIEJvWO4po89WBZ9ALBFN3ghvxsJJtnbB1lLC1TP8vuvNdEDaMRugIZbC4anhhl7DVwHeNiLNNaZXyvG7EGOg9aAbyoAzlJT9BCYE29ELDQq0Z/EtuU34ifhgfK+enJ9KUHvpDOnj9D0dXUAThdAkxaxYtnYKCTJiZ2pNvvvJvg6O00y06UGKqZHrSGOnhu4R5iWyJAejtpfKNY0Sdl1CIeFTAx7WbelNkquuzuhAPo9+zKfNCwnl6W7qTIrGBV31AE+/d6y5Yt6djJUYatj+fzAfZMTk6mc+fOsTHAbmSAHKDVYn7045mmDPUmWqEPU+T1HA94Gh3p4MkGqMKYyE54dcK7gdiZaeT10s//5A+nf/Ebv52ePjGZmoPjabm/AweMl6AT00DwzRQB/ONaDukz/dL7ybXX7c4wXlksAzWWV4+4a9j0HRrsMB6McuyUGECKgECMEWNbvQ9CT+HVc3guwnvMT9oPPYqVwYBHjpFgDiXjfUT7XgsemuybqqkHqm0FKINcPPfoxzweZNMLgGTsNzJ+YF+66vqbU3tsM+8BwC683tqMbag2tJRn9NszvTU5F2Iso111M+ulPDD6LMlcxzHKDpRRXj3kfaUvpLv5GmcLsqkXvrj+8cBdKwH0oGf74XGGXFvEOhPoMuaceuDyQeeGMlH+c8RVs2/KShm4FFYwzk0dTAKZSjWXEezLchOslY71PCIkIQXzfI9ZF/3PfNIv+qs8TJ71KDTPsVcNou+MmfM7eHOuw0eJG5frUjC48Wc1nxGw7+yYPjyOmHnRSm5nrT3GfIV2pQ3HUUKavqdyGVWde/rHziuVvlblIG4p5b/WD1mpknlIKO6kGffS2NDnUjb6ThnBb5MyjPLc24aP7JubU3iNmOJsE+bFLqvodC6ntNBfeI7+8zLQy7Zqo8VZz7ERwHj+0lR1movnpbV+5L7G76vnFahvagl88yRQtOybR7GmVEuglkAtgVoCtQRqCdQS+A6UgAZAGAHrvGsFeoTZyDd69/z03BRBhaexd5cNar6EsYfhtYrBRlWMACwFjZsIcK1BBMBQPMqCvq4dUNOU1lMgDCHqhGEHsFAMNY2HMOiqs9flXn40noMSy+MmicV0+MSZNL5tN+AYRjBgTUMDEkSDxMZ7mr1h5I1MTc8eGBweO/DGe+7BsowyGjx+D2r3fEekNVspuA2DHv5d62bY8Nbs1l0H0n/z3/5K39Jy353EZPs+rLGbWH7WJG7WAvJexttGoyzGVZmaimwFLZW9S5j0lijGtUa7IEwxzCzjEWPNuSTlLNggvVLXc6aZaXtd2vPaVMquebtgSaovWuWeSztQBVTIPFtPvcnlvMup0LeNJ554ND351KOUY5MHqknHQy8eepluvPn1aRAvsdBXwAmBAL3spJm9RTJ/3sdyLIhIX8BLD8ZBYvG1ASGGCLKvB5lLLfUiM1/QY9hll0MDxAgDtMCxzzx5dsmlHkF6Z42OjOEdRpB48k3yLY9TU1MBmrQCpOsPbyE9LfUSU0568Zjmq6WWs+zMaDD/Ii/nnqnBHO0X4OnOpW0j7fSLP/3jaaLDGBiPDJQ7vMhizCisXGg/ZBoyYIzlS+GRIlw6GxUsAKw9d3o2XVgErMMfLTXwMnOeVUCXHl1l3lvPvnkEAOuw4l1XPKjsa3kOFBVtl77lZ9nTyms9xyIv3h3ZU60EjTf+4MIy74OlRjozz0yY2JmuvuXOdPWNd6TmKO+FPmLDtQERAccEVJXzRj2Mca10U569j01BqrzyfOO5lMvA/bqeKr+QIQUCCIOG8dYE6ou3W2xqYp/os2OqvpWxtY2ojy4pmwsXLoS8rGv/5dtrduaNuVPkJz/W894yXqurAmVgdZFKn73ZeF3uoxA/1njYcK03rrRtmxL8yyBeqVP6XM7mS6ck2/PYmDaWNV8AvMjY++iDFyTzN9Io9+qT15aN8utNrrVf2rVcoRUXG36UMr6PXljGevlY589760hS0M96uf38BwDBvI10fFYlLtfer4NcD3O4e3QIp+JxQy9KtfpcS+BbL4Hnz9BvfXt1C7UEagnUEqglUEuglkAtgW+aBDKEsIHc12RsePa8Sz+BvsFnkJ/mGGfFKAj4iPtNmydW8cQSCVsVTPAjvyRBBr1s+vEC02jQzwDzIYwGDas+vG3Ck0gPBI74a3plLBk7Sm+kyjCIs6aj8cP0lsjFWLIGMOAhkIadmM5PzqavPv5MGt28Pe3afyB1hlmlgrFetQ85zE7tJvP6253uav8e8IS9v/M7vzf893/qZ4NfemBvn2+MfG1O1c2/Rm5FGN+kcxlO/WfysYHwOsdYaFj/jVb3wJXXp1/757/eR+ioe4jF9H3sMfrqBTxOqthZfRi2OJtkEEVKekG4y6P4V8bAaCUsVL0jNKApw/1667n/jlM51IFyXc6FS5eweRi3THDLccnlHWvvHUv0hr5sHH86BLIgXdvLhnh4qjiYcsPZZYYa6/ZHXTC5e2UbPdKr6sjxI+kL93+eJYgXAlgRqVjq5hhNPTwML7vq6jSB91YToNddJAUB1+ihvd632UlSKLEAhvKlzIbxANs0PpxGiBFm3CrBswH62cJAbnMMAZZtHhtO48Qk67A0chPXQ+H9lefLfOURtASfg8Qwy4BDlo39EDybnp6m/8yBCiDroPcd+BwA7HAnRT2OTMpzlqWWxiOL3S1ZhljyY6dKwCTHb8hx6C2kvVsm0n/5Mz+extjjdXV+KvUtL8Zz5ejSNneMDYHqNcShN1WhJwDQQyC95kg6jYfWMyfYdZMdIW3BsY/xDZBODxnHT1J4vqkv8OlSSe/tLzM43gFlOV3MWZB3PaTkpQCViAhwyGXaCxnopq7jFF50lPNacGx6oZeOTS2n8yvDafe1t6fLbrknbd13Weob3AQwxjixkYFLXjMCAy/que84xtkYY/lAH5VG9V4L3VcFEUED3XI+lIDsysQ+57J5XtiH/4+9dw2y7Lru+3bf7nv7Pd0z0/N+D4DBiyBAiCRESCTFUBKpF0WKpEJRIiWWothlV77kW1Ip27JlO7FZLsexw0SRVKVyPqQqUSVO8iFRpSqJZEsyIZKhI5oCCRDA4DGDwTz6/bh9uzu/31pnd1/AUlIlYUCocvbM6XPOPnuvvfbaa58+699rrx3JycSha636Gkqk5iBidbd61NpP6ziWxhNLoDgIUy+TYKoAmXJRbrZpPb3Njhw5Aj1kCr8uWzX5h4fKl8tyQ3dhwXZiOTOEfS5w5tlUY2eFSJQA72Pjjykf5+a+PHiPW8V5GXOFNgWB5Mcj+tbMRetEOzwf06tRGfOuEbiVl/22eZ7XCXIFQ4x06I9n9YSfetXF/KN8AFGwJzBWwTHbr6kZvuA78mnbvnj4e6X2J34PNbKpvMYYovfRloC87y1lwpFlqAAPHvJhnh6rlkRS0c89dBzXuv12QjY+pX1/L+olp4esbU3gvjre7U0BrguQMVVSpzy3qZXAd0MCTq02tRJoJdBKoJVAK4FWAq0E/v8sAb/E/SbSEvaoX+YDwANi3/vB3ilnzl0Ye9+T3zezuLQyzbI2Ylhr+GBQYvkAbkSdMHw0DqtBwnX1JrP8gXGZxpDlu3ikuHucxoYHVkOAJZWWwInsVcOBm0ju4vfNZ55nUeF0ufTAO0qP3QYFPrSTMl4PUE/YTB3sk13ije/oSHNiuz84xa6F0x/90Y9BJ4ye2t+G8tvxZEcODMBmhJoxw9Ld666fvfxg+eW/+8WJ7d3OR9b7O5/Fm+hDW/3BkS0QQWWHDHocEV7Ee+VbDTzP3ntUL66Qv0Y0R1xTpwIG1jd5rtdhdDbAQKVf63mu16EzDmmTpGmq51rWc+SHSnqVOiCgpnFeDfAsh2wEdACWNMC3+hvlqaf+ZXn5lRejrPzQd9QyvcROnDpdLl6+h50jJ6O/gjH9LYGX9FZSHgILBgrPa4AGgSo8wCYAWSZYNtyrwKI6Swr6nAVwBQMEIwywf/jQbJQ3mP/EhLu/Am5QZxuwwzbU7yr/6WZHQoPrBy/wE3KFP+nHZgeUn4LvqemJkGk19jdZvrlJ0HqBwwCvEUkjQgAQPeZYYkvcq72t1fLIvRfKZz7+kbKzeie8yHaICegwxKgySWyHBkVGot2QLZxvsMOmXmTbeJAtE/T+hdsb5Q5eZMYlixYEr5h09if5llYje+oF6CF6Qf987vJqj9Qh7o1RCA2TxQKEAVBwaaL9ql5nW/TDoPzrAGPrO93YnfLWFoDRhQfKI09+uJy855EyMnsUN1d2eDQOnChnk6qs671tZ/s5hubXvHquZQU48g8BQ+BSU7/q7RtpOW7uegr74UXmtWCvMrBsj/h1dSkkmSk3GrSeycD7gmSm1PUE3bxeWFgIGiGnprw0fVZ5t7+mkD2DrE5UcGy4rGWqLnkePix3kBoAh3lpmcrnQf18t9c6lQ+fv/E6gvRDu7YrrXptn+yH88hEj+LePMvUPsZDfki78lNp1PaG6Vq+5tc6tXx9Vs/D5YbzYplnIxN3rq3vzFq+8sar83V/CLIdj1pOYBNtwKN3dJIxfp0HGeUoFsmm29RK4C2TQHwkvGWttQ21Emgl0EqglUArgVYCrQTeFhJI46thhc/4sI0PrKBcxrZ3/uI95VOf+unyrne+q5w8cWx+d33pxI0Xnz8yhjtKF7BBWIy/7ANEYe1hPLr00b/07xHrRzAsDT6ACYw07Rzj9YziyRJGlcsgKWF5vTjC+NTowEjyuUaGuxVG0jANbwyMZAynlZW18q3nXiosEiuPPvZEOXycjcBc+sXOf2moa6RjUGEYQ5k/2LNXIcbh7s72OGDfYQztaY0Xd+hja7xsg5rBkHdNs82DodPr5DaU/xZfJn+YugizdDfuf/R95W/8nS9O315a/rH1/tanMVHfhyxO4WVDz5F6GmUdjbkYI2QZ3iTIGxMsAA17UJewmaf8NeItx4ikgjAOGq6CBJEATzXAI486KAH0EpgRcNGoDbCFeupH0KSi9EVk0oMDXhgnVcj8MBl5bPmyzUEb6ocp6sGLlE0HQAy1GMcRYk6pc9/64z8q//fXv1pWllymiPcawJYy6G/0Aa0Olcff/T3l7Llz1O/RxQHx6ZJ2DcAvQGUKzxA8h7r0V6BYWQRIplGs3sKvKKzL/JSB4Id5epPYBZV+Z2ynHMLjbHRULyh3bmW5ocgt/dMLyPEQoFPnxw263uU5j/UWsqzJ/rObArIEuENCsTshixunplnmbOD6/fbZzZA+OnQRgJ4LPc76AErGk2NXV6gxt3bWy0c/+GS5+sr18r/+3lfxbjvO8kRGmWWSTMhs1zkJ3Whf/VEd6M+2W23Cx2hvunznteVy7dyRcrK7XaZGKQuQ1WViBfAnEyTlbrKPjr+8muW7IOY4oKYxz+yv4JibbkT8OfoOrJ3y4tp81gdHfWN4bRGbbQ28d4Mlnocu3FsevO8d5ciJM3i4Yd4Re60uFQ2dsV3HRaVEfjoejdk/bsmGZupeRQljXHnAkKMf9sdxEgzSm80xth/pqaU8BQH1vLTN+u6Kdmkt9ICzdY2XJz3pxpg2Mkn6yqeXOk1h34vSWl5ejF0svY7Yjkx5aY+zXHRubi740rtMXangn7rqXK/zzfeo77uITyefyDveCc1y5QpOH3CrXNBh5wH/d5H3DrwKvDJ6vlGDN7rVyKWCYhQmBYDE8LtE1Rh43ttHU7Qbcx8+IoO2nOvMml2X/FI23yMpOWUlOC3o7D/fJ8lvPpeEqeqZ9XeplGOa/Jj3+jK+e+S5eY/FU/vclCfbKsrcs/MZEcYRciFP2XY5Yq5bCKViC8qgEb/nqBMLUXnme44SjAE9CP5pOcYgQGAiknV67BLr5IxJkzKy3gH/eY0StamVwF2WQAuQ3WUBt+RbCbQSaCXQSqCVQCuBt6UE/BDHbhE/CWt9F8gLGxJvEAJc87U/9rkv/OLM3/jrfxNAaaSsraxNLt++/cDqWv8SX/YLLN/rTgE64Eam4aoTGYZLAl8BZmBA+UFvwOK0MtPQGMFjxqU7tNUYb9Y3K8GTMD4wOsIucGklBoo2g4aR5pSBnldWV8pzV6/jNbJVHiHG0MLp83j6QFfjE+NDo17jw6SBo2GGYWeKvM3t/vz01OyR06fP5LP+tv2uj6PM2/wHndWi7ICedAdXHnl3+ZW/9w/P3F7Z/CGWmn2SOEffv7W9Na/RbEIWutCFvD3XANkaeMrJuEcm7zUq67UGd4wHY+zZ55zi2jHLlIayz3WKcZxMGvdYqVEn6yWNSo+H0MFwply2m15DLpFE9cJTyAFBqyQa41jHNPIbfrJf8I6eadzqPSag8NRTXy43b90IHbSe5QQnRtm98KFH3lmuXHmAWFRTtO0Sz07ZAvQIvikbdDCcwYIw3KlDXug3GfI6zTJH1dokOJa0BccEb7LPW4A+sVEAfFp/Ql3m2O4DLyCoxeWl4M2NEwTLpBEyxGPMs6CESwjpGfUw5qFd8900oM+ySIGvsptgid5jyklvI5NytN007JO2M0gjvgPQ4SYFYwB2P/tTP8YGAbfK1569gSrNANixSQb1BKNoMJematxDb3/sUD29yDp4Zy2urZaX72yWh+fxICMeoHUIQQ6Ix3jQXNVB52CVU/RTVihrkH3zAxRF38ilnp5kbiiB5xjvIvVKtaQY+BtjRbH+Xrf02Y9i4sjpcvbCfWX+1IWyhyfpgFVq8h5ej/SDXTpCHgI0yX/cxrXiEDSriVtFGMmyJmUoHzkXBHAYK+5lxiIVJLNNJBvt1brWF5QSrFEW0rGvke/8IKlPLq/Ug8xrk+XyTFnourwy5ZEAWFIoscOqMciUsXStX5ftCeTKe+XFZ/IbnmP0svKBZkW9BItSRrZfebW+LHuf1+gO/bS8+TF2XNR2LJf9EAS1wexjgFvQqnS8j0FtJB6gYdOGZfwnTXnOfqVsIg+heq5tRXnq1BQ80bb1aj/rswM+6/uw8ltL+M4xZRs1t56VqTSlU/nynHJVLim72vY+nw179T5aqP2VlfHRHn+0iSD90mjKcYrfz0G38tCeWwncbQm0ANndlnBLv5VAK4FWAq0EWgm0EviuSWD4gzyZaCz7vNEW5eN+VOQAA3ekPPHeJ8ov/uJfmv2Rn/jYicmJqTMvv/zyYWi4NG+aGEAPsgHivZjegC+boyx52usRC8mv+F63hy26A+DkLpRBNAxbmwnPCgwqjYua5CuNCAwUrSBACmySNG7D+Enjy7/wexi/TOBidWW1XMOgv7G6We5/9L3lzD0PlF2WexmYXyPWpikYRoz0palxOUL/TJriUJwh7/j65uaRwVb/NpWE1niqbDTHrXV3Uxph/98Nvb7c/thxIXzT3XrvBz9S/tqv/L2L128t/SyedZ8g+8rOXn+6Lqu0L6QRZRNGPj0VrND7xDGoY2Ke4xbGHvnbAdQkf7WMQI7go/WUlWWNLSfAZNLDSaM4nsd4W8ayWoAOC/QRbR5CKIwpkvaIBHhjXQ9pe+BDlI8YXw1y21Uf5DX4pXLKSIO8EG9spXzlqd8v3/jGN8rG2noGthcE459jf+XKfeV7Hn83O0ceQ+WSVizbg7LyMdbVGGBFxKNCX/UM0pAXeDOO0hTB9nucw0gmf5f2wwhXLjAgDXn02CSeljzaH+U7irfiIfqwxjLFLTyjOtv9Moq63V5apN42nmPqaPZ3FH01ZpbgR5U/UoSPBNP0ohGsmWTJ5mCQ8resIKDLD3GtinhbPdTEwPnSkD+6Ac9QUu60eWR6unzhZz5Rnv6Pv0QVdsYE5NqFrxBmTAXKIacAROibHkihR/DZd0Dw2Hvm5Zvl3cePlsNT7GRJ++OA4CET6g3wbnMJqfd62clp8sI1fTBu1h6eWAO2xwzdY5zcQAGXJbzFqEMfdwDzXI7KYtcIwr9VCLI/jdfapQfKuXsfAiPEi05WGOc9dEOwKXB4+tsRRLRNGnYsajJgvuOiZ0/oEpyJ51hPADk8KRm/l+jbCy+8UM5fuliOspyxgsnqskmeTS7/NM9xNiVt9SNu417vNcfN/nc6Lt1VL4gpV9+Z1msO9Uq5q5tLSytlQMw6RrCw3h0dQG8Z1/m5IzHGMQ8om2Bvzp0x9CdAQvLDkxbdl6fgC9nWpY22aF49B5gHjxFDi1yGM+RChdAjsmL8hckihhv3IYlGtlUeyjI8g4O2tTLVuaOHVU0xlxgmdazOF2Vl1WF6itpDfmu+Hm4V1K/0PEsn3vuUreVDJ5tCyiraohxNhayG6zNC6ED8rohyFgqQj97qeWjyjzVe+vtNXY5+NP1NmfIM+Qr+GQjTPxw5ZVJU+f5S13pshUvq8X5NDzLmp2WkIY+mg+tsu74n4mH7o5XAmyyBFiB7kwXakmsl0EqglUArgVYCrQTePhKoH9gNR6x0HAXHAObASuYmPMZYttTpTU5Of/GLX5z91Cd/+sjm5vbZpeW1S4uL6xcxBxawlib4vu8RRPrkndWlC4AgU2vE/5qdJLA0Rv2+MYD1sv9hr2HGB75GQ3o1aEjhWSKQRSGNvzActM241uCR1/DOIAtzM/JymYxGhUvQRsqrr90pL9+4XU4Tb+vc/e9gZ7pxQBTrGvxYCOTAsyDa1kRJI8mWKq/TGCOnV1dXT9HmKtTT1YrHlnl7pugHY2dnOphZo4PHn/zQ6C//3b9/6dXbyz/FDoI/w8q3h13GBjg2oM8iNVpeAY7ZJ+Uh8KOsPTT201hPGcUYIAIBEPMFCToY/NbTQGav0hCNxq+Wf8iV8p4jT6OuyWcgIq+2VYEBy5rq8s5oh5GL5bh4B1ne9oK2dHmmx5X0gz90RD3JoYKvGF9G3ecY2Xfu3C5P/eEflOWlO9kHKiZo12HHv9nyvexaeerUuZQBm0mEjtCmKQGy7dLbxvAlYPruLvmJrwRtg//bDzVZsMIUOtvwa1+61JEraQUIw7V8m4w1NbZh/xKIYyoEoHLr1q0AiVxehhUdQNYUSzK7LIdUDs4JoSUDuwt6DLcp0GW78hWyhS2XeQrUrK2zAHlkqowT30+gxWXO8hUeafAzYnv99XLl0kL5t77/PeWf/W+/H8syyyhzijYZ8f32YTDmrEscYQiPT54Dpu2NTZYbS0vl5sp2OTsBgAjgw2ap0d+OmwM4nvCzYz/Uo6HkvR5Y0R+XpnYtE9ALdZjL6NxgG3CM9nbY5GGdcdnqTJT50/eU0/c9UrqHjpYN2ve9YAxDkxsKCDpAKfrpWMmD98rH/pter0vNPe3R5f0+v/LKK+VL/+Q/L7du3SkPPPJwIf5ieeyxx2KjhAHyTJAs9YARl2r0Rfr2KfoOyGI/a7uOuXzU5/5BwTF1DM23jjz73CRIeOfOnbh3KXDk86zL+B49fiw2l1C+plo/aDQgi+QERX0Hu7uqKduofEdW/Mg2k7eam+0xDsaGoy/OJfnLseN9MjQPhvvl9T4/MGCb3lcd8L5eZ73UDfOcxwJOVQb2IWk17xxY8D6Tc598uUIutc7B8yyl/GteLRf1Gpl4Xes2hOOUdbKNmm+52h/Pw9c7vDNNtQ2vfW7KJcUxByFb+Y+y/KWi02WOqsQwkv1reIqCfxJvQbT90UrgLkigBcjuglBbkq0EWgm0Emgl0EqglcB3VwLNx/UBE833eBgK/PUcdAQDpZR3vfs95S//5b9y8nOf+/SV5eX+lVev3zhHKJSzBDM/TaD7k3z+z+K90cXYxyoYneBLfrbfH3QMBu5yru3u+MjoOIZnY9AZl8m0J5CA8aHXjUljUoPbYnqMaTQEnFWNAYprfGns+dd9l4J575Ivy/bX1xIcu36jLJy6UB5595Nld3yG5VZ67WjASE2j0o5W4wxbA4NFa4SWwyQRSAAzGqeO8blOUfRFyrOdXzBJheBfTsiAp/jpLrokBwAAIABJREFUj+yX0N2bkQ7ovoFatZuaAsPlkAcdQ6Ajvf57fuCHyl/75b/7MJ5jP0MXP072FXcs3ML7B48dHJ4QCqBCn6V31ZjVEB9Dti7RC1AFo9zkdQfXmZAVY6ZeCIZFHChu1CUPJRwADnX0qAKXoFx+SgveRHlKhcFIWc8eQT+MXoAAxBgDwXgJkmoMuwHEHvcCGwIjjhFQQNxbOPQkOB36IUgDb2lkA/bRB71/vvLUH5TvPPs0HknrpdsEvBdgm5yZLR94/4fK5cv3ymHQdFmihqcx7YwrFR5Yel8N2ImScECCeHtjgBHooP0PLzB4FHBQzQTAQufoR/UeU9OUqoCQeg7eE3NjrFnyaHsVGPB6nSWKt29eZ1MBvN0APfSccefWCZYKHj58ONrVeyo2KaXtHbyaTPJjfduzHWUsn/0m4P365gayJZ5Z48Xmcz1q7EOAENDYJb6b8xTtLz/6g+8vv/MH7Pgp8GOcMpZ37jl3AXBohNLKW3BMfUDQxiGLcRsryxuD8uxLN8vlQ8fKHDHRBnubeKfJm0sit6NN25ZfGJV9yOTSyioL3xVeC8LEONAeoC86Rp+Jy7W8wfgAhl185D1l/sw9RF/rlrUt4hHyXvB90RvfC286d/kcAUgSYPmT5qoxsWIMYj7Lo4dySL2j2XivreGpKs8PPvBA+fKXv1wuXroUgN1v/dZvlQ9/+MPlyOF52hWBTtCxLqc1VpfLx52q6j7CCM85uhLnnAvoEp5tu4D+4d2FTGJMnFP8M1lXPt3J9ObNmwlwqmesqpasMcQM0C89y+m9qbzti3Vrv+xvxsrz9e1cA4CUQNOGZ6Rst5vUvN+QB51AlvLNuHO9HWOWxfTc8tCrtKZom/bVlsqHu1YGeGsuk8G5J38CoSbIRtu244VLg+2Pt7LpEe9s6qvn0oU6RyZBVH81VY80yaJGIUdpI4mULYSsa154REb73iQwaTdCr+03KX6f+VjGqCcdfydl+/BEu+GpiHztcf52oYi/P3jfkBP8Kh/rjDC28qj87ZN9jCSvuG73t7ZH0QGe2Fp91OhmLRsPpdHUbcq1p1YCb7YEWoDszZZoS6+VQCuBVgKtBFoJtBL4rkvgDR/RYVkAeu1iTLqdIxhLd/o//dI/OfpjP/Jjp1kp+eALV2+9i4/5BwHHTrDM5jDG/yw0pvkUHxOowmjf3elglo73IJHLUwwA35mb5INdI8Cg5U23wwII6yIy0qjIj/owjjAf0gzRcEhjIT3FNPTTuMSaCLMt1oBCZR1A7qVr18sAD5Irj76bnStnC3Y5hgkGIsCPXjbaDbYShhA30a7GCUkDVHBAuewNdidGxsZOs4TtNA8nqLysKUWb9iAZDc7fLj80bbHIOkRv3x3deezJD479h3/97zx0a3n908ApP03/LxuriaV1G3R1FH+dnkCoS/BM9r0ut7L/joGyGD6n0YpskIBGtyZmBVOMk4VZG/LFxgu56ucT8mUsTdaJdpB3tMFZmpap5yjID+89qnEfxjzdS6BM/rKOXk/SynYYGK4z6WWStOXTIYNcWVy6Xb721S+XzfXVoK8NPGbAdni8dOFyuXjxMjSgDa/GvjK5HFG+Q17MC41xr43/ZcB+k0uoerQXS6nsP/zZbQ32AIKtbzmYEIzbN4p5nrypVj4HTFpdDdoCB9Qu2wBZS3i9GcusN443JmxJZxJwrwdQ5VylweSxGc+klXnKRKlkwPeUqfwLVlpXGQrCwCKyyDp1rHZxnHQp5x47fi7MTZV7z58uT/3rq4DSbnSA3DXokZPeWQNjtEV/Yj7ty2wED9JtZHptca0sbh0rJ6fpA0q0ya6Y46hRj+fyE8AE9etYCj4p9zqmLptlZCK2Gr4+6C4jS/lNkCUgu1Im58vDLKk+deWd5cbKJkHr2ViBNlx+yf8yur5B/0pZnZkqR4jL5W6htAbgQj/UefqeuiRdhy/1VH6CJ/JCB+BJvgQbL1y4UJ4+dqzMQu/SpUvEPXwhAKt/9X99vTz8jofK8ePHHYocd8fBdhg767sRSdCjneGkR6Rj7egLVAuUwRo6mTqfPMqb4Fm3bGyu7+9gWWWnDrv89ujRowHime+cMdl+zgnfpRwxl+hvqmDz3KHM8vLqtYdtDx8BPDV5Lnt1jJDSvpxsbzhlv9OjuNL0LE8BNNFrOIxryGabDYHabp0vApb+njGofdaHX/RKOUnzjcn6th8Hulv1TcAyZUJ1+0LFypM03kjL+rX8cBuWi7r88Hm+I/Pae5cC1xRlact836cm38W1Lfkw1T4zFzosPR2b1NWT7kZDWYCOsjizGZtax3ObWgncTQk0ans3m2hptxJoJdBKoJVAK4FWAq0EvqsS4BNbC6xbHnj48fKrv/FPZzc37rzr5z772U9s7+z+PH/A/jnsiB/vD3a/l/P9GGCn+Gg/xAf82I5GsrYJn/t4c3VG+YbXkNcIY1v6MJY0FqpnRjUu9o0BrFENgfhDPHaBnhSWiXKcsYLwUNBLgTYwwDQzrAu/UcZd7NyJ8KVrN8rtte3ywOPvK4dOnC8bfYxuGBOogXoY1J5NGqamaDeNC/oORMRjPVd2dgdE8t45gdfRSTJwOdEOiTYlEEQ0YdKMkZKZGDjBXd7ftZ9vaFh7CSHBE9b0SHfvkSc/VP72F//R5eW1zc/udUZ/dm907LKeNpt9gjjh0EKfNcuQXXQDLxxAkOqVoYHYHIJfgJ0Bgjl+jAjX3bi3uTqO1dAM45QldeENgqw03gV8hpN0gpbjCqCkx4V0HE/r1brWEVLyCJub9qxnebsr2BP3SDxAKJTScbNWnhOQsw/BK0vztgZb5atffapcvfo8fWT8sUxH2DTCJWrGG3uUXVjn5g6zNK0HQMXOiKAq6pj/BNEEd8eIc7evM8h0x90KkSr4awAm8mRfcqmZmsoD54f6TX70dR+44yn59klQhC4EWHV78U65BSA2jqxdsrm0fAvvMeJLMUaCCBPTEwGOGbhdEESAS30OnaYt2wm6tO6180Yg0DbMj9YEYJC7IFR4YVkGwz8AG86W06C3rCBYh2OK18NjD95XdjZWyi6gjIAg5GOTjB3AQstBgIkKsOWZ8bAN+etOzpSXb68Akm2U5a0Bnl2DiL+G9CjOODfAhe3qmdOHhrrj/K18mc/mGQA5PTYJYHko8dRW9FLdAYAjxuBD735fuf+x99DWNMHpD7Fclg0F4BEvV9hKGRnz7cZrt8rTzz5Xnnn+almFD+aMkqIvOXa+L5SbKTwY6YN8xTJe3lX8ESH0otsDN0dnTwGSnbt8mWWqvfLke99T5limOzd/CIBuFTo59kEMni0v+GYb9qsmAVP77HioT7YnD+5gqgyjffJMPo+XGRPBMq++9hr6uhHzmLiPTCv0Bt3Qe+zEiRPBq41KJ+YeBIz9VQHwqrPSSn7tO8repCoLeYgkosMRQC/j7JJtU7xrGz0MftVp+mmqsq20PDvXfQd5rZ5V+uHB1rTluymUN9o44EmajoM8SNu6xrHzXSE972tbwQv3KTbOdI/Syb/IKZUyrlqOOVJVsqF/0s74YQf0lGO0z9k2/KVBy5nXvC/0ru0x3noN1hRl4j2VIJ356kCtG95p0AmaSS+I9vn9tj3o09re+OyhGZR/x9dN9IPCXKkf2b4029RK4K2QwOtn41vRYttGK4FWAq0EWgm0Emgl0ErgrZEAX9aYKR2cwLBN3//BH5j43//P37n8sU98+iMvX1v95O3FFXY8HP1xAkx/P3F+LvE9P4NR28NbgPBh+F2ELY2ZogMWphtGV/w1exRgwg/93UGG7tIWdLmbhkc1hve7J0CgAdMc5msPaRBbVu+k8H7RRCCvpjDew+rZxTNopby2tEbcsfvLqXvuL2va5xiKmDWNJcFpiL68mYbOZhiLy+Br8FrG8RA6iYF56oMf/shUWF4USPMqrRfrvw2S36mI1XVV3c3zVx4p/8k/+M9OL6/1fwRE5WP05JKgB8a3nmPY3wNWU7HfYNN/lzFpKHs/bCibV+81COthOeVY63t2TDXKLe9RDfFq+FX6tU6OYQI0lg3PtcawHW4nnjV8xqkB07Q5pWW/hsubV/WjAhMa2y7hdWnoyupi+erX/rD0tzejXizNoy8dlkpevnRvOX36dPAviOLSSMEKdWF6ZrJMAUoJRgk82EfbsW2fOwAhq0YZKg8Cc7XPAhoHwEfquh5IlX/PJgEg4425ZG58nCXOADsvv/hSADyWF1BKIIBdL/GAmiAOmSl0thmX2r5nD3moz6MwPxwvPeCMhwToHSCZYIDJOm4QYLKeANeusmBzgvvvvYTRz6RjXgNPBNAStEX3SPQ4foIuZn8ByWKJIDJ2yeMLN+6UVUCJAeAGSHqAFDWmoO0ocw95cBmlZ8dZACCeoa8CXgHqkdcHIOkDyk4fPlEuPfhI6TdgR+gvIp2eYtyI66YM3FzB5PJU2V1cXSvfeuaZ8uJLryAD+uq7hPoCuzFu1Knj5/vH66rLjpf38n723Ply731Xwpvw6tWrZQevtWee/uOyeOt28G45y9exSDAjQY0AlQQikbPPTfY3grv794qopw4nuGW5Wla61nGJpd5bXquH6ojg7sKRIyzD7aGGB/2oPCRPyAId1RNLkLb2ybnj85q8rvfW90geKMNkjD7As3nVHSrGFICz1qs0htt4I/1apubLU82r7fpMOCrPNN/wluOSfFunztHa34P6jtuBnls2+IZgLSuPppofN/ywbH3mteUP+pN1oix6Wee6z+XFVHnwXO+lY6rnmh+Z/Eg5h7xH19fXJy9dujR19OSp+mq12MFA1UrtuZXAWyCBIY1/C1prm2gl0EqglUArgVYCrQRaCbypEvBT5k/7nMFCYk0Kn/p7n/7Zz4/99//T/3w/u6B9cnNn+5e2dsonVje2H1/f2Dy91d/uDbAqMUEEj/jZ4YRxwW14aPAEIwUHLzyMuuN7Hbxf/LiPGGQYvtUACCMhvBn0jEgDKp9Bm0/96jGhcWR9n2lspLdBAjV6wuzsErcIA9JrAumXO3iQjU0fKg8++h5WGGIAw1sE/cZLQY+0MHYwco1HIw8aSdIOg0cgg3VGxjYDSMG2i+D1wACdozNzR4/9F7/2G9O/+Ff+PSwcxOhWY39K8rHHXUu2/G+2zsDuKsy90+zW96Vf+81jK2vrP0nJT9K/SxqsAiEAHGPIYCSXBNJf5KKd5vI5Dbh6yLuy8V5AJuN26TuWGpSxijQyPcjDAIxxjHrQRWout8t8vFSinTRcBUo0vn0Wsqf9Wk7JpTeJ7ee4OO558KzpeK2rfshjNTrTmNZ4Fyhw6Wh6k0V/oDMA0Pn6V/6wfOeZb4NACEbYhvmDcuLkyfLY49+D7vWKy1DVFWPWCVTMHpoux1imdvTIXJkhKP8EXkLy56HXj/zsG7w0Zl13K/QcB/3yeeXbmGU1NpHPzR+WvW2uri2XV6+/wm6sd9gd8TkAnKuUY4j1YkO3x3sAdjPTGWoOAUEmjvACRPNN0tUrRsnh48M8FXGGb2Rhu86fmLzwlkBZ1sPj0OxI8uK8s3z1Ujt/7lQsi9wdbLKkcit2TjQYvPJgevFuEGkCHMMniMnEfQI/8a7oTpdvv3KzvLas19coQCVAGbKyOdvwveJyVPXS9nJsd9DBlHkFzsz3OZ6t6BveY0B1lx96BLTHeZ/6o+fYOMDYVG+U5ZQzZZ5llZMAjmgMZSgFZhExwbh49bXF8vS3ny83bq0AlCEx5kTKWwAQevwQlHE5YR+ZmGL8obWKh6x8Pf7443iNzRMsf6k89dRT5bd/+7fL4uIyaomeUFtHJZN8b2712Rxhg/4P8Awytl0u4aWBmGfO0Zh7yBVp0FaCUL56Rr1GYB4uv3Sc19iJ1T8obOMxqzy7bIIAhwH4jk8IXAsY5aBWPVSGoiz7cyi4S72Jd220K9MMiv5dMa+yE/bdtMMc848YecAT13p8pUdijrtls/zBPRn7Ou8mLflOSDnbL5P6EF5djK90k07TPs8r3QTzGuFajmfGWqvx1vwLTsYBpI5ebzwzqZfJ1zCt/N0QBfhR29BLLTzmGEnfK77TlB1/ZWB8ncO2ynuP95HyjUnmr1WuBfNrqu3JQ/BBZ9X5Ot8cZ/WOHjgPcF4MwsjXeTwyir5PnTl7YepffuXrox/9yZ/KiugkY6Oj4+tSbet1me1NK4E3UQKv9w1/Ewm3pFoJtBJoJdBKoJVAK4FWAt8lCeQn9cgolkunfPwzPzPxX/7arz+4vr71UTCCj20Pdt+9tbMzto0BIOSAwYJJq3nd2B58gQMyYBnkUh0/+PU6GRcE0WsBY5VNL8vyymKADphEjeHgKY0HvQyME6WBqaFGU3FoF2gghbFhg83Xvx/9tlM//r3WU+IOwbJvrayVh977wTJGoPV+GB0Y9hp31gnXEIEE2oOWRpMGdDX6whijPZcdkewjUBKmzUhnCgbn4X3K4O2//o//EeQa48aSb4+kFLH5R8pPffozICi9J9jA8ifo+PuIrTMG+LGFvMC1cBmij8quHnpd2PcAGsj3Wl0wv4I2XgsPhEFHf4flX7uvQ5GxoAKwbJafBTwlPer6z6Tcc+wcf0C0MMJzfB0Px2b4sI7ljZXFidJp3NJak5/lLWeqOlONUu+7LFETPNtYXSlf/9pTbEiwftAf9NBA5g+/89EyOzcnVZkpWxsAOHgBuURPUKyL984YwO8oy+ZM/f52gEpeC5IpEw/b2yFEnYaz3ArMikuEvLnOYOHJu2DWKGCLU6jK1BhYGt/zAC0ulROwvfHqdZbqrUcwfueJccfYKRY2x8r0NCCZ8wd0xH5E3EDoRfNy0PAVS9FGBJwcj8wP7ywsc2WrzAXD+gA1PUDROk7ybZ+cp4ILI3i3HZqfKvfde0/5+revUk7+E/RRX6RBBRpQJspSXgTgiP3lnO5OltduvVpeW90ux9nddrKjp94W7Tr3Uk4H7wIAHEjYviDuoNlIQGBjsItnGXJSBtv0YXwGAGzhGPHG4EdvQcbRPkyNTwSguLaxmYATfVvbWAe036IutPFEE/yw/2vkvfjStbK0NFXOnjlVpidzebAyzB09KccyXfu3Rz+VjXxNTfFeox2T3pjuYLlAcH5BrwsX8LZjQwDl4jzaYjno7cVFPL7WAsSa1DORsfRZtgOoh4ciE5I66Q2m7In/GPRtE+HGtfKWbzda8A8E/iHC+wR+2ZACOicBfs2TL+WYoHb2t8t4GNsMrgMEVfdSbw7acr7J13Dy3uWz6j2ii3er79XQE9qQiHSMNxnv36ay9SrP9kO+nP/qn2m4HZ971LnFw9eVifrkZLl8f0imgvbmm/K573/1XtmkHKqMlK3tptxsI/my7nCq9Mwbvh6+N18ZmPRqC6/J7Frk+cPn6kLMk/3c5sK5wpz5E/gJ9snv8Ktucn1ja7o3MTP+8U98qvwv/8P/KNXgqbZdyQ7Ls+a151YCb6YEWoDszZRmS6uVQCuBVgKtBFoJtBJ4iyWQH+5vaJRPcqKrYNt8+vOfL1/6r3713Pra1o/yDf9xdut7EC+HMXc71IDEWMN6cA/IBK0wBghihcEx2NFBojHmNGr0WsEQwhA1ePIYgbzH8GbQ2Ksf7OklhDGBsQIAhdGQRodGiyCEni1hzlBfQ8J2PGtcVeMk/qJPZwb8NX9lbbO8enu5HDt9sZw8f0/ZZhe7XcAi4xppo8Md9dL40V5xqV3sPOgSMKxyDYvqTQY7toFBgnmNUdkj1tFoZ2ySm/F1lm/OEJ9qbYVg6dITHJD8W5le32DgVkAwdNBP1bHpC5fve2Jldf1HGZNH2EV0TE8O5Wd/6BllAG2QpfajRwImabjaDcw6SqTBpaEeO1lqOFPdoPUa6gGeSM0DIpAPOYYiUN/d7CyjwUppxpOC/peGIIsN2xZ5srR/r/DJqEa8ZRjxALO8DkMaoupHelqoJdmXjvHTGFcVR2vSMdUDx6bUG5fWvfDCC8Qeu2oB/ssZ+oMO3HvlvnLflQdKj+WTgoOCUZuAG8Ya03tsYhJvHvQEsUUfJlnWOJidiWv75CGoo46ry8NJ4NA+KiN5qs/tc3IgTfvAXGLQAm+mwjGCvguwLAKmeBxhqZxgWB8wJLyLJth5kvhXC5QTMJN2yJeG1GnHzRTzMTy6aE3+4cXlyoJjgmmCdIyUzEV9+dIrSMWq45J0NN6pL6AEnSfe867y9W89xyM2JsDbqc9OkYiBO+c02cqBt0V2njGALwFHl3Wyc0Z59pXXysXD54hphtcNBLfhx/huXbydHBj7YzImV8qt3+QlX4OIycTmCYz5YG+8HDt+okQ8MBp3p9FUsQQbpDvHMtRNUP/wKGP81gE4Hef1LXbYJX/AIY82u7yyzrLLF8qJ40fLiYV59EdgxTlBP+hklKOdkLd9JambKf9ujIfjV99Z+RzQlTZv3Vks16+9hsfXRoBLU9OzxAhjV0/AWQGqPYRM96FH/Cq835xz0TD9lL7vJOelgFo8BwxcYYfTPrLdH38BQpg1OP/CwlHAL8fUeQ/vgrLQFMjm5c+Y5lxvuhE0YszsLEfm226Oh1MsdCq5DKDsABxj3IJHeUWvqIxfYcw1gUz1yXZNLhelt0FLbzVKxbhHLEFoKIPoTyNn72sKvZQ/xtX3uO9ix1j9jPrwygJyePE9xAN7ATPGBPT95bsj4gMGK+qTJbIF26zt2p5jbXu+wuKdz7X3vj+CD6kHgZSj7Tjn3aDDMayAIMMWMnQZ7J8UqP/g95CAu/xkauZ19ALZApDtTuB/OsnfPHJnkGjf32rZvrzXVPnzfji/Pm/PrQT+vBJoAbI/rwTb+q0EWgm0Emgl0EqglcDbRQJ+f/MljdcREMTY+GT55V/+W8cAAJ7EWP4hjNLvYdnPCEY0Ky1H9jD+jWCtpUEljAWNJT7+uQiDxKUshnyPz/qwUiSNgTeB5013PD7OAWuChEaGX/tD3/GSJSPrJ3iTxqbtaGSEwcLZD/6a57XG/t5gpNxmaeXW7mh55P6HsLAnMQQxCOFTu6Xu0JiN5E9pNvZQZGQb0IMpjb1sB8lgSOrB0GdZy1R3/NDMzCHsnojTpu13YIkME39rrxEOFuLoGOsnu+VTv/BLF+9/8OEfW90cfJQxO5XApsDNzrh90bjWsBZ4sY/VeBPcMSl75eszywkwCQ5YLoxsnodHD2U1AjNf04yR5wcR6ZAhwBRgnQa5S4/cOdSRdTGuYxL/lZzeEuiCsu9gsNqmqfJVDbrIhweN2ppi/LjJ8UrgwGeW1bTO8czhsT/2z+Ppb34Tz7D1MKr1uNomb5T4VO987NHwznLp4uLyEt5O2xHjaprlupOTE2HIB9AF80rKOGTLeADZjnRtQ0BC+SXfAC30rQsoIPiVqqK3U/Isn9bhYfDsfYCCtIT0AxQRDNOL7IWrz5fl5cUItm4ftyk7znx1bGb0mjp6JJZZSjyAQcoIKqrHAtHyE+CNvDkfaNeYYybjmA1cpsw/+yL/HhGUnjGvKfoUdQGUPaM/JwFexvE+0mtwC88r9lqMtjT09a5yoC0b/Xc+CjiSsUsw/JHedATqv832sodnpEHbNoaO9GKcc0xDrvBvqjorUT1G0ciyAe+dEZbE0p2FYycZG98Vznnalhz0sv8InjLyq1ePgN40BdfwENvYnMRjjDHHk81Xl3HWBHcEk66++EpZ5tmRI/PlCJ6DHQBTwZwAOChsG0op2kg2vYt7foRMQ3bkDkImXJB4nwRYZ+D1DTYIEDg7Q3uzs9OxsYl1RgAOhZCMJuZYswtCjF0sfWSsuvTF8XQO3mZXVmPWJSAEI/YfOQnSzUxNRz1laZ6Aj96QAmMu1VRHGLJIPCJBlHKWNclL8MN9vQ7dVVeh+TpwLO5Tt3xBmgKUg8fU8cxU1wJEatqRjuNS6Vu2XieVnNvZbvJkPr2ALnJiEJTDPogpOMwLScAR0vu0rC9dk7LzXl5MyYN8ZluW85nnKgvLVd6a7pnVlInL1/Ur+tnQd9n5Hnpb2690rDVMP/oIcYbH/GhGOszLYJznvc3NncmZWd5C/H4NJcym9zUwbytfw5zWJ+25lcCbI4EWIHtz5NhSaSXQSqCVQCuBVgKtBL77EsAq4P/ICLH3R8s7H3/X4dOnTzy5tt7/wX5/536WcIxss5wpvKoAEgRHOPFtH6GcwWPS8Ii/etOXiCETHhQuu8l6BsHWaBFooS7LmsBwMB71uRr1r+xaNYIkjSz8C30ksv3re3qIZbwX6ejtYpKGQI9l4KjcIcbPTY7TF+8vhxZOYXASlwijaQ9D3BrVIKnGDjlBx4Y1oIxNYz8tpz2iucSyRJmIcgI9PJ3s7+0c6e/uzC8vsr0g9rOAHq1Y2i5U7qPOW/Mj+ANbGGNVzvjIo9/3obmf/OTPvYvxexJb7JIgAp5CfQwqC47t4Pljsp8aozoVaWCalI2AUTW4vRdE8DDeWLaEJx/ddDmsSbkpf2ECzThC2IXRvYNcNPKSsgAC4x+eHBqx5mZ9DXStO3mIHeLQB9vtoFt60QjSyKvSFYTgNvmjvGBKGpIJ5AmexH0zJnqxSFePsj343epvlBvXXinPPf8sNbOu5ZFVuffes+WBBx9mVWovlt1FcH54U29nZln6Bs8CTqEb6iZgjzrocwP/B6CEAJTfAJryHHnUE0gJ8JizAJj9RXJxVozqfBca0lQuzo2IT8bD2ekZ4mX1yrN//Ef0XTAD7xfouGR5imc9gGeHwB03nR/yFyCbg0Gyf/LimMpP5iUALP/mx2y0DIejUWMf2WNBotpv6wqs0ACHINFeOTI3C994lxrIH4+wsOVjOviDcvAsYOelZ8dDYG6LPkxPzJSbeD29urxVjo/hpdkDqLQNZGqS3wRmBSCzH6IgQR6SVcYuG133+QjedIeOoCsE/Lcl+Ax9gJbvCoETGQm91tWIMuZ0x6YBkCbKoelAbA5pAAAgAElEQVTxsglY5xLFDd5TAajihaaQfL8sLa+WG5NT5cjC4TJPv3t4uTVipkx6tjIhoHigW3HDj2zbtgCNkYO7j87OzQQ4W/rs7skfDlxuefXFl8JDcP7wXHigOfdMzqQRAJ94myEkx8335hbvZ/nUK+5bTz8Ty9iVm3h5D4/dLvUvsLOmSXDSJKjmMMY8bt5vdezVId+HNTmHQo5qJY2GLmXjFElPLPU36tMvweYsJ4NIu6n/+sBY9EbQmOfOa3rGP3VL+o6PWpBAYLwzKCkPtqE2On4CX+b5Kok4YHFtGXTM+em73zlGX6znuIRcbNTfGTxCJSiTtKN8Q58SUcb5EZ5u0DIWnRM15Zb8SioY99Qogm8yqnHvQ8goZ34E72Sqj4Jk0b7XlT+r0X5snZxVY97tx8mUZlB2GqFju3vjSGgS78eeILqJIvyHUCQ616ZWAm+RBFqA7C0SdNtMK4FWAq0EWgm0EmglcNcl4Gc8q1FG+bN0p/z8F/6do1ubO+/Z2Sbm2Nb2UQ1ZDRYMi24YGRTWEPDwI13wJT/gBxhjeI5gQFguPvTDa0ajVQOBZUAssRSAcjmTdqp5Ec+H5zJRDQy/8b3e0XqJfI0lC2WbLg2S6AhtacCYiJFWbtxeIubQZLl434ME/cY0Euzi0MDLFrKNMFCaPtiuKfiljSyb9xpOJoybKKaRs72zM43ReWxldW0Bqa1QJNGmKPld+eF3KcIYJcR5d/fw8TOH/v4/+McfuLW8+qOMzYN6zdl97S77UcfQMdFI3gZstF8ajtiAIQevh1Ma0wBWlPPQSDRZTlNsBIOf7T7DgI8H/Mg2s5zytp6mLVs2AO7gacVdDIv1G4RIo9Zyjn200xCr9wIrVUe81vitzwRe6nXAOXQGMnISfFaQQZ154fnvlDW8w3ysN096JI2WJ598Ek+bExFPbMWg6S495PkRgIopljFW3tCSIT1JUESQTCDZMuFJQ7uoJEsGs591ToRcNI5JQY9z6B7MOiYCBLYpFKnHleVnZ2fLlXvvLX/09T/kWb+swrsbCMyzUUAuHU1QzOV2ykB6ghzS89ppFLLQc4V7x80xcXml5wDzmjEKD6Vkzp+kamwz7I2M98fT5ZAsSzwKyDNFwPtVGhGo2DUofwMYRoB+eIkJz7tEEMJYalBjV1kAU+brRhkvVwmMfw+eWfP6sOExZQljoKkayiDBreTfvgX/PHfZIbvpolO8A/AcPXzmNHHRjgKGuvyWeip10zenifU8h+x5FEtI1Wn/w/soMcJ8j03QH3cN1YNwc93dPZVZgqAuD3355Wvl1VdfLYfo++HDhwGyxtmwAfkjk4j/FiBR8ptt5hjYbtBqxmiePvsHgHU879ZZaqlzkMcSu/AaB216mrhkxDRzbK0bfDvGzjbO0hIc20IWArPPvfA8SzbX4pnzQG9GwZMTJ45HWQgkmIRg3XBD8UjTJBAZc9HZqRto4P08J7/2IQqGTmTf1B31XT5StyA49Nzy8ulRx83mEiTOZ75eaxlpcAOtfAeZ77hEfjaOQqReh8cbz9xcIfC0kEkDnnFtvw7oyW/WUwMqz/5xI14Ekacssr0QCQUF8mEhkjLwvWOSr/RSax5GXuZHOZ4H8Ne8KwN0hKg8Kat6SKvKtvbRs96BvlFrMs93DO8kcE98cOEFkHWc0ASHVlfWp53rboizN2BnVhm2s21qJfAWSqAFyN5CYbdNtRJoJdBKoJVAK4FWAndVAvH97/f0pz7zufKDH/nxuZXljTOYXyc3twZdDCBtICwxvtn5aI8gZYAufuBXbysBE32Twj+JonqRYQnkAWENtTGWBml8e2xvN4aghDG+9BrS6sE3Jg0a7Wn+CRJkSmOwGid6dblcD0sgDDx3fru9vFaWN3bKhSvvKL3pw2ULrzEBOGzN/eUsGhke0gmzxmdQCQORDI0OAQr7ZtK4xBAKUCmNSL2pcNcpuwtT05NHcQV5WbePxjNEkh6SjBRtcLWf0eT/WU9/Cj243B0dGZvYPnXhgfKlX/+nFzDgfxyvh48C9s0Zg4lEgc4YBjRdUqZpPIZ3DMwJVoVRh5W5B8gTAIYKwTgYH0hwSQNPA60ahhKtBq89jOGuoAgSHsVi2434YKkz1quGoLJURYzBkwk5qweNoSxdy2skjsKT1x6m+sxrwZEE2gBIGOgwLMlDoSJfMKbWc0xHMSDX2eHv+vVr7By4DrCAhyHAgjJ6/Iknygc+8APQGSkrG6sBMrgUWF4P4yk0xVLKXgAFeMdgtwZ/DLe6pKdXHMgnDFfaMnB/f4ylhNSnFyEf66R3HRJzXujlppyhYT/sYuRHXx0YcukDEijn8ABaOH6s3L75Wujn3sggls2dOH4yADSDuwtkHiTp5tg6lyJOklY0yTYc+2qkh0bQZreZ3+EFShkgD5Y5Wof6ypR57m0nAE6AFuaX/Ts6N1UW5ufK0k08Q8PbCYqCYYyvc2PPOGCUc4bvOSFN2v7wIxQ4wi6cz756uzx4vFsO4ykncKPXmTEP3WnSpJhCVMgiZSYJgAYA3gDw4X3AstjjZy+X0fEpli6iM7CBCOP5NmNddcHlnfY9l4IH+aAZY+p4ocfqnro/3usDUBFnDnn16YegqWMcBzQWAeXv3FqMstOAZAJZ44CXvufUVcgFPbigfd9vtnfQB/VrcqoBv3huO/IsfWWuN9tge7OMrLF0lXee5aUtgFT7Yx3zr7GBw7Vr6Dbeb75zjfvoDqcnTpyIAP3RP/64oLed13EgxQSBmnv5CzVhvNjp1DK1v/Qg+Wr0aCCIRVnHA27jDxr+gUHZVvr21ne1/+RxFNn6+8Ln6S0qp7RNu/5uEQxz3kY9aauF8ZoIpsimbDzlChqmkAt65K6RAfJF3/T2QgeRodTsg16XwSvtOw7my5e/JOTN90b8jqMF9Tbed5xjQwpp7rdMPQmQZBVtaHjJcXXGC+hKU7Im3xPxezLmhO1nfZ8EkSgTReP3Tnjlcmsf/SOVtIzTiW7iCAvMv8NGEswP+nV4sLN1ePHO8iTLmTegRyedXK9PVVYH7b7+eXvXSuDPK4EWIPvzSrCt30qglUArgVYCrQRaCbxNJODCLy2D0fJzn/95YxpNDja359itckbPhgxyLRBAoqQf2C6x8sz/ABh8FAYG5bu99O7QINZww7WI4PYYRoATuoNoH2/hkaFRGzHJikt+NIrSkJFO0m68YJo2fa7xpKGjWYP5F65b0tN77NbiShmbOlSOnrlYdljm5a52wEFhK1R68imdNxo6jb0XfbBs9KUpi7URVlg1EjmPY5sc4/ECBtT4oL+3Ll1SYwrlzVvwU760snCe6Wzv4T/205/9/KnZ+aM/sLa6/n6M3sN9dsnDHtukDJgHAonua8RxhZFosr/2zfhqgkWOmTISCBAoUBYa+hqLlg358dxkPe9rvhQtLxBQjeTgMErnMw0/JWodU5TnMmWe9Gt+pVvb3C+DCtQ8OfE6wQjbppuNAa7xW8vV8Xv11WvlxvVXGmM1gd65w0fLxz/xyQA3lgA79MCxvO0LOgl+5dLQlAcPEmAZkofywd1I1tGvnANe43EYNKQ3hv7nkPnkIIU8mvEwN/uZMhKk7eLR5A6EegK9/PKL4eF2/vzF8sB9V8rly/dE/DF5DW9OxlHPFb2QHD8NeCWtHCzjIS+Oj6nm2UfnRc2v5dWHHjLwbB/DOwxgrMEwmF+DMsFujmeOL5TnXnuR+oJHADbojN5UezsAU5YXGLDNmCUwiJ4g4YLaEox/trzGuFxbXC8XFybL7Dj6M9iAfxcTAjLAc7xLGn7lPz2d4B++7d8WW9VuA0zNLZxsdq1liJFBAHTUVy+EcUzqhf2uKeKIcaP3Gw94zzB+yt2xH5sozHhirRkrDI/CSXafxKtMOQkky9cuoPL2Vr/cWjdAfj90yzh7XbwOjyMXgU3B39qmsrUPjrOeaspS2drfASCc9B3DPjHJLOc72PZGiXsmjU6zQ2WOUXowCszdvn2bTRyWYgn6BJsPuCGK8+Ls6dOxIYHlQ7dQOJfGCoS6bLDqm2cBKc+WVZNtLzwi4YPMpg9DusSQxpJs+qD+xdhE3dStoA0p6SXwRb/DKyvHJPN95u8Y2zzQVQS5f+9FlZ/X0lWVKgjObUN3mIYlSfDu75voC+fU0UYXYrzzWfVU83dX6m++34Z5rONmK1SNVJ/n3UGeV4Kc8W7g2nKx26f8MMCKtKboGwQt47Vnk9chw6agtLb7W4R0TJB2Y2Pj8HZ/4xI7iV6gyHc4+pUG18FmUzVo1ev23ErgzZZAC5C92RJt6bUSaCXQSqCVQCuBVgLfNQlommCdxYc4uwyOs2RpeotdDzfdtZK1NsICYRjwvZ0xx/S0AqDCANWQ2yZ+05gx/jHy42Meg1mjNlMaAn7Y91i+pIGwiXfNFkZfLEHDGyLAGgy2+mGfngQYTRoKEJGSO5JpM1RjQcPBJgzC/dqdlbK0PijniR81NXeMIP0Yaxi7Yg7V2PBshh4FIxF7iFuMDI2hauxrsNug95YXfLM9yrGK0OUtm4A7u9290d4RDJ+juEwQ6IhCmSqr9T743r/5f73Q1BtOQ5bTUPZ+S5knooFMxvBgc/y6x578/g/8xNLi8sc7YxPnB4ydhjU9HsW47giY6I1kn00avS4J7APqDBgPkwCZhji7osW9ctBbxXGpBhs1969ziSzyGfSRlfRTbhBHbvCG5giSaPgKUOR+pEE6aHQBIur4mKusazue03tMT6U0GsOzSV64N0VZ2g2dEIjh2T49FZOWBQhcLqZHx81bd4jR9M2yvgoABrgRsfUAWD77uc+XKw88WG7iDbS4vBK6gwJDS7dJQDLBHuQVOgRV5WRSurU9AZvRLiCigAlPRvBgFCzRo0UQRZ0Llqgnn2GMW597adgHgQbp1H7EQ7oRu0saxJ0dWmkl4km9852PlXsuXS5H2dHSMXLcNhg3ASV3EA3vvCCuFFIutS3nIAzYgWhXcMz6ehx1AVrIhFcAPVxCYwdAxjPkqDyQhSn6AEFXO09A675L58v/8ZWnC+5WICZk8mx3Vz1q5Eaf6Wi0KU3nXbZDEUCoQXeqfPuVm+XSidkyhycWpcukbQGwS8vq8Q5q6ikz3yEu791EzzaYA9NHT5TeocN4suKlir7v7DXgO/2t8lUWOtl4X8czl3wWkGSe0tAobfrcmeL9GCCSXlB6lPVZluoSzPA8jCWqyJ55NL47HnmTzAXfM4JAOpvq2ZfjK8AsUKM89ISkLRrYpR3Hbxtg0bOTSNBP+uMAhS6DFTBzbjlGwbNg3/5Y6OmWnovPfvs7bDwhHp7zzZ1XDZt14eI5liGic8rOBC3nozqoe5Za6DOaJaHr9Lm+J8yBy4M8dEv+qQAgJoDHOyVAUYfXvtl29lOdl7ZLIE1uBJDeXpbhUAbBa3NPufqOiue+10ghNy8UGEkPOJMydJT09qOUncr3eYwcPNBPl14nGJWAkuCYiR4f9LF5n0gnvfSiSPyQj5oCPBTco8/RlnJyLtkQSTIhO/KG6ylbWbZYyAqVjvdxyKv5Hcd1zAkJ1fymbeec40G2Dzu+ijZY2pyevrtzO/3th2nvmxR4jRZuQUgaIXTyeTU7LlFZAm1qJXBXJJCz9a6Qbom2Emgl0EqglUArgVYCrQTeYgnEl/0o3gzshFVKDxtiQrOJb/LGKCP2O8ZNGI0a1c23th/tGm0CAQbEdye2/bhGGAnWD2MC+iMaPxhXGg781Ts++KW3/+GuMUQFn+/nwUwYbk25aiDargawwMM6nht3ljfK9PxCOXHm8j44lmaH9A/oSbsedrQaDp6lWZ8Nt28X4IEQW7lsiDZZdbZ3GI+NwxipWrRQirpaSWkpSfyuJ4S61+nuheXVK7/4V//9e+bnFn6Ybrx/c7M/1d8mKL+RwYgdhzE2av887JvjFQZ+A4jZN5dl1cNy5pmUid4puXTp9UYWwwK9NNpDdjyuMqzdd/zMq23X+yr7Wr6e63PvvVa+9bqWqePjWRM7zkNjW8tbP8qiW57XV5bxsLnDboVrjQx2yrsef2/5yA//CF5jG7EbZYCiAA6uK15cXIy2a188S0f6ccZSjbbEcYLf5Nl2Q36h0o3cwyDP+tatkvRagMP6psqzZw/zBbCuvfxKefbZb8dYnDp1qpw5c6YcOnQol79aBhqCMS5J1PNJUEKAudL0XHVA4LPKrT53jKVhm55rvuc6dvIiv/bNvPCeAph0qdzl82cbMDRqMNfxHlUfnBKUzYMM+97wtQv4A0pS9thtdmxqvry6ulOuLW8SbF/vUPLh0rK2JThS+bLdPui6cdiMM+jSysVNYsWdOAPYNo4HGfpLU1ar9SvPzID9pXbOAWmZLFcP24vxE/gB/HJTi9zYAo4oJ/Ckp6yedbFxAwBGyM18/ggwDsDnWEzPMB6Tk/tLlC0j2FFBRtutMvUc3lDozHA5+2x8M+OheR2bZXAeBQT0PsaczRr0ejQmWsgKunqsCeweJsbZaeKPRVvm005c2x4v8tqWZ+cyUnudHCxb5eL7u14rH4fRe7Up85O21/an8iKN7B/PmYtey59tekC2oeOYMWgNPeuZLC9Nl2/aWsaJtFwCnf5C8g83f1qSZgB5AWTBa0O/8lT5FQAzJX/1fEDX/Pq8vvdq3Urr4LmcOg455l5H3+JdlLLx3uc1eV/p1fyQT+QnbzwnxB3+2ICpTfmZlZWVh3YGuw8eO3tuRnBMUJBOCJChrslHbaM9txK4WxI40OS71UJLt5VAK4FWAq0EWgm0EmglcJck4Gd+fur7SeMHNd/lGJzbLOnZGeD6wh/n/Qs3Di0aE4QN4prMgX+6tiJ/uecDPAwbl8wNiDXl7oB6nG0BkullUQ1PDYdqCPixv7q6Gh48/c31MOAF0CiRxpqxcbCW9BDQGDNVoyFu8HJz2aQ8mzY2ttlZDo8fllSevvxAGZ2aITi3u9dhNMOwIEc1ODKmUAIAggMe1eChVHgzWLYaFPkMAwbeMKQDIPMZYABbRe4c2lhbmt3pb4BCpCFFRaokz8HcXfhxQD/GjdHpbY90Jjsf+cnPnPj4xz/72Ora5v3s9NfdJLg3O/A5NLu585/GbIJgGtKbgJkbLL/cIB6Xx9rKOp4nCZop7z5gmYcAyziG2HC35EHD2kPvqvDywxA3+Sy8OQREm0oxfsooPBTT00UPG8dcfbBcHY96L40YL+hkDC+N/SEQifHSOK5t0mroatRXN6nn4ZI0lxma9Ba7fesWAe6X8fjpE09qs5w6c6587he+wNjjgQTQKqgyyTJGdV/ATCDXBNZESl3yCmGGnoQ+UEcb12a7GOmxbI3e+UxvlQQSsnyALvaWPsdzvU/g0/wqO3fbFMAyRQwsdknc2Fgv/+L3fpdxWgpvveXVlTKBp5aeZeGhBwOCIXo2hdy4lh897xwjhZPDISBiHbpAOwJvyrUH0GJ9ZR1eeoxtTY5fHUvBZpP3zu896Ao37O1slUuXz5VJlvW5pDJlpfed7XBv0H7BF18o0HPoBCyKc5V28c8s43MLZa30yneuL5YbK+gmuNUO7VQwiR7RUgJzwQT96ENjlYm+vAXoOzpRTp67VEYAzWxG/uTdAyFHs9YLfeTdIsDmu8Qj8hiv1OcEfHP8sr0cR8dSWaBTsN5Dbl3kRUzCMs4Y9cbHyoRx6ojBNskulxMck1PTeOSxA6zjAr8CWsoulntCA9dPNCW9g+TNZ+qwSz0t6+F4OkaepS0wsr8rMNc9gE09j1544UUA3duh2xPwZDmPixcvxhLc8MClnCNb59n+fGnkYqwtghkyVglcyZNejXQ7wSnHk8P3pR5v6oNexPlcnUbwzbxUfvYj3u9Nv2r/YnksvNiOY2O+SxH9LVPH23xpeCD51HXKWVawVBry4hLkzEOS0oz2rcsV7LjsM+XtmfFWnxGCJRPkYm5QR5DX53EwL713oG3bPPlw3OMPPuTWsqOMTfOrSnFF8pmyrXI20/HzvVffB771TPFOsF3K12R9Uz3Lp9cpG65UG1zXxnpjvN8HE2xffJbxuPgbv/lfH378e7+PitCqk7USbc+tBO6yBA40+C431JJvJdBKoJVAK4FWAq0EWgm82RLQSPIw8WmeF/zs6pExwH3DBUJ8kIcBgmFg0og0z6MmP9z9wHdJ3jYGqUapXhkHRqleJhhS2qgYBGMYiv5h2+fG7Dmgh0GDMaMREiUxFjQGqsdZZPIj6WY5A6gTHr8sr/XL7LGTEXtom+BguxhdmLhRxfLStM3Kt+c0utIgsqD3Yag015UveYAGt9lp+4f31RjB3afPnTs3e8/D72A9GfQ05qLukHAk/CanRj7CNdieo1hxvcHJM5fn/oP/6G99AHF8GJmcHhArSQ8x+jPOWHTk2SVa7hwq4BNeYuzQ6H31oLHvXjuOlrG+SQNPI13DXJCoEUM881r51hhAysryJvnUPqt5GqOW93EYjViani1nfj5LQ7neByF+NCSjbM3zbLlGHpHtfSxR5Fyfy19t24D8eFoACK5GnybwuvnMz362nDx7jmWVqxHHbgRj12WpeOCV6y9fD3nYB2l7NmWfATuafPPkw/7U/lree8tqwAdYyziIWilrj0rHspWG1/UIoKsBSZbu3Cq//8//RSypcnwEmR3HAFAaPmxPpCJ29BvmBcVUBo5MNdIFLqIc+XoGVjoCKsP9lab8yGs96tIweZaeQJvHqWOHyyk8lQQbBMYEEnaRuTiDwAAxkhTU/hEOLoAirgHcRld2OujY7ALLLO+U60t4ke0w91C6uvmC7dm/6Cdgq0urB8zrPZZnvra6VeaOnSnTc0eIv4WHGO2lDubZOZDgTY7VQV8aAIzZaz8dl6pTlhmmUfMtV8c5wDB2rtT7Tk8x5TcDMGasuJkZdvaMjRP4e0MIIXoQNKVt3LMK5Kl3mSowFS9MhQhnyE3vOcBe2zbJizxUPtTXZ559trDULp7Lh+M9NT1RLqDfAkchN/JqnXpvBemqA55rn7P/zbtyaPx9nwuO+VywyVTrVBmZJy3bsL1673m43XjAD8vWtofl7nVNXmfvm3dIUyfAeh5I13eRSVrDKeYcvytqPM3hcbacdbN+vqOG61Za9VzLDff1jeXrM8/ONYFsr+uhPta+1X5Lw+vhe8tHv4f6w/NY7s8Ys8dEZ3eUcUP3jnbGevf2d3Ye+vwvfGE+fnETiwySKE+k1wukyWxPrQTeTAn4zmlTK4FWAq0EWgm0Emgl0ErgL7wE+Gy3D/EBrdFNAhHKj3lv/EiPpTjYOcYlwryPv6qH8eYzPt41fgfEIdMzyYD5GgBx6H1AGYGBODBs1zHmVgApIoYKRk/YQBi6HYP4h1kHsIBRoQEZRhseFqYwKCzMYcyzjc1BubO+WXZYnnX20n1lbHIWLwQMaupVQ0RvmGqgaV4J+Bl/ySOND+81SmwjDVD7oxEU9TC09bKxLODRHiDSHm0DOu1M3HPf/VP/7X/3zya+8Jf+KkLaN8q4+rN8JmoIDh/2+E9NNkA4HwK3X7q//Opv/jfHVtY3PsTy1h9gl70ja5ubu8SPY0h2OivLa507d+6UWwTvXgIE2mRzhA0OgbA+XmaOWX9zu6wBlm0KcgKSNeBagAVVDq5e0nvC++Sz4a2OK3oR+oB8lfG+LB37SOiJ/aOcQFvSyXPIWaDEg1Tl71lwiQVF4S3imI00R8TQoqx161jblLsqaiMzkvuHdNTfAAQ38QijoEb+D/3QR4jldSnA2xW86IzZtUX/lcHVF14qV69ebWSA95q8ieA2/NumRnY1XgOARU/Rtuhb5cn+SC8BmjR2nQeWt8ywkWxZ80wGuVfO6t4EoPVXnvrD8torLxGo/3Q5Dhj8yiuvBH994k3Z35AD4oViHNZ1qBw359A+AAZyZR7TC8AF2i4HhH54JrFkcNylmZahgOMtqCQv0q9jJn/VOUX+o694500xfS+eOw3AvkV5ZU47lB1xGSW7XsZrxv4xHlSKeuqw4LIwpnHDutNHyuL2aPnXL9wo15bWyjr66Vgn/+iCoJhAIwkYDg8zlsKOTlJnr5y+9wHmP3HAAG8sU3mLTQUa4ERefbellBhDaMfBWDr+dUzCqwyeTFUfcy4IpOQ7pXpzKRs9ycaR8wwg2dTkBEvV8SJDtj1i0sE1YF7zlg2K6ERtK3YDTT2QvsBW6CuD5PgF+JwXYoPBn3pnst06trfwjHz55Wu8E/HKVb7W4ZifPVTOnj0d9axTx9BpGx5Tjc76LMbR93vwlJsPmKd7lJ5ezasX2ZHFTdzLC2WqrCv9mA++U3kWnmvSp0KAWYLjSMUhSUArwbbooIxEoiwF7KOpGb64DjrUFYS1D+5IWue4BaIObRh3MMdTwNQnCcj7uyr6Cm/q58GGMxCN3lmW3wsAarEclXIVpAzZ8sz+mhS1R3KZOu0z5WBZZnlcBx+hB+ivOidF+DP5TD7iYNJwG3V9FjSQQZVvbRfGWMY7EUCsYCy/puh39/ztW4vvOnJk4QFespN47EKYP6L4KkzykmxTK4G7JgEVrU2tBFoJtBJoJdBKoJVAK4G/mBKoX+Rwj3mx3wc9HkisTMSCI/nx7sd+NSjiQx8DIM4WwKDYISi1H+4apQar1pukGqjhOYIdEF4nfKd39FDDQLC8wMH+B/9QW9XIctfL4fY0FqIeS3rYRCB2qhuMjJf542eJP3YsjOWwyjHm6vLM4H1o/YsGdm2z9mEY6PCZxpvJ57Xv2e7O3vrmhiCZBSbxRpjtjo1P/+THfooAzC7rFFJ4KxLtYPjsYsB95ue+0Jk+NP8OgMnHgcQWAMcAuza3ATp39IpaWloaERDTw8SllSt4Hin3CtrUcbKvAmMBjg2Niwa7sZaUfY7LgfFnXk0+G76v+Z7DOqOsxS1T5eq1h7Kt1/VsPa9NlvcIsKCpUw3nzJdOAprWcXmumwdUANFbUNEAACAASURBVMGzbbiRgDGvpDM3O13Onz9fjhxeCE+sAUZzH3BXPX31xk3AhpcBK8YDsBCEMO33Ed3zuh7yYIq2ybc9n5mvbnm2iEa6IIdJuSeodmBSWF95V76999BLy+WVdKKcOH6q3HvvFfgn9lh4Y6bXk/RMlSe9wwLkgo8eYEvIjnkX9OCvC0IS4Ir9wLr3sI7tJxild1KO+Rv7ErJsxszuHOgQweDPnglQwLhcukftspQ1+9HoB/3xjYP+0mZ6k7r0NgLRI/u9cUDu8bny8p2NcmttpyyubfG+cPxSB5SlXq7hwQS/zv+bK5tlm+WVC6fOsbRbPCDhCtv1/WQSENO7MAG/fH+Zn2AuF1E2dU3wovZRoMwkLeVgqmcDx2ffEjAzX69C47/1euqg9VJvoyI/pFvlpfdVrIHmHMn3liAsqbZv87Zhv7M/eR/XDVBnu9evXy+3bt6IejFnkZFebQsLR8KTTXrqlXRMlW+vrV9pe28Zy5uv/ubOqObFLwbOjkXyNFzW69fTrzwnrZTHQV+Geai6avs1VXqeoyyse67zy+sefYo8PLToRVzvy26IH3mPfMWLnGuyrvTtq6nKorZjntf1qPfD/azXw3S8tk6lV8tU3fJZpeW5Pq9nea1tmlf7XPlsyvH3A5fd4sRM4v0+y/t74djC8YUP/fBHp/cYp9pOFGh/tBK4yxI4mFl3uaGWfCuBVgKtBFoJtBJoJdBK4E2XgEZCGAqajkb64WOaw3hUmBwDAAbC46SBb9suc4odKzEwNOw16epHvM81ro0x5LGzjVHLUh8Nwbocy7PGZgePivAUo8W1WMqHBxgxigzoHUcYiBhU2nECbYJp2BIRHJoLaeAdhRcaIE8hBtD0XDlz8V56gDcJBoHPaWrfgJNPd5/zrCdbgmEJ2Gk0afUZd0lDwv5WT4VqnDRxbgizpdfRgA0KB8RjcwnjYGJ0rzM71unOYZzixIARNTaKpaVFLOG7kvz+pKHOgF3/trvzC1NPvPd9T1y9+tL3A4qdWVxeK3qLCYotLa2MuAxPIGx1fS3AMUGyCowJhDk+W5z1HMud3gSRHD+AS57paaQ3kWNrSq8mZZsGZZWRz8wL+TUCFBioyXLG6emoI1ybGCa6QR7dGT7q81o3PACVrWKNsxUP5KvB+DqjUa+VBjiwvF4+Lm9S12Ps0bURdjZcWrxVrj7/XJmbm4M3d4Dci51V3eXy+vUbIsSxo6N1BKiq0S3gaz+RRvBU+bQtxRR9gSdBJvvoMkBpKGsPS+hhqU7XA3WKJF11S53TIBbocOndt575dvnWH3+zjOKVZKwrPUaOH10g8PrJMjs9E/237i5zR171Ohun3wIkglw+UwbGyBK8EQtQTD6LGGcAbcbT8lo5Rz7PYlke96HSnO1z9j35VSYCizEf0Bn+lwWWWbKdBV6JbMLBM4Y3nu+x7LcJHB7jIwN6ifr2kabHjjIB2Bk7dKQs9UfKq8vb5aVrt9FP3iPISK8/tSU2AaH8Ku+B1cFYef76cjl5/t4yNc+mstJDP+A+xiwBCvWVZjkEdnx/RUJPqndo6BBjGDv5ArA6TjUJbA6/6+Q1ikLQcVe2jr1LIMcAk8ea+F/SDB2QJ2QVXrbML+OO2Z98NwoQcw3YbRvqyjaH8SB97nJp2+jqBdiMpXSzDWKP0ReB76effjrq+ix0Hv1RTwSBBbhDl6AT/aRjsXQdGQnohYcXw6t3prxU8EteQu7ofACSvliRrP3XIy694hjDRscr7ZgLVXy+yLlWrzL2ne9Y6ZinvDnihvxGFzJD2SbQbDlqU+Hgnm6i69JMgFf1rHoUOsXk8k88NlXl7NlJl79i0AMacr4i1v15Y1vxrpFv9EiaJjdmGEE4Pg9d8HE+irysl3O91ql5nn3/yI86rIylUZPPR3kXqixRlgepowmy13KerTdM37htpmZ5L7/IRwdLK6vlb/7K3x5/6NHHxvSojl+AijCLRvn2RyuBuyGBOu3vBu2WZiuBVgKtBFoJtBJoJdBK4C2XgB/eGjGkba43/VjX2CIJEMWDagRpWnhtHUEUwS0NBg0OLKa43tMYBBTQMAmjAoO4gzG+hyEuOOBOgta3rsaYZd549rnJMMoe2hUaa30IbGBUHsFrZGScoOqNUVvbsp5eRJ6lKR9hXGgg2Tip0q7X1eDZz0cWyXcu61IExrDxgGaPjQjmMDwX1tc35wV7sC8xgTBEMmUjzc2bdPL7E0uK026H4PK/dJTg8t8LqPXeW4uL88bX2gI4BPzqLq2sdJYJRr+4vETcraWIK6YcHEUBBq+HjwTO+oKjaQQSO8rA4BrWjnMauDne6oUy8vC6HvYxZZeGpHUirykfN/ywfAevoNAXDdzmMN8UzyMv24nMJl+jtbYXXhVV2uicdASIKj2BHo1lj+yD47dVFu/cBki8FaCG/BqvygD9d5ZWyo0bN/aX/tquhqeB123LdrN/laM8mxdxhigjMKZnl6mWDw8cumaAd+VseQ/lr36Z5NG8eh91qeP5y1/+cllZusOop3Gsl+cD999fTp44EeWrjtY+Wsck8OH4KQfzfK78YgfG8BQbkhWPBGEsU/sqV0mrGUf4q3Q8e8jzgPlgN8T/jh4+EsCqehQ8QJOCMpPAuPmCAS4zbdqSRgUEtgESerNHy9put3z7hVfDQ+y126ux/HIEnq3nkltQKSZbtyxuFeKPbZcH3vk9AHE2leAX0g3+lI30a/L95BG60/Do9XCyvJ5c2XfBk+x38pn9trzPlaUyU8655DIByOE263X1FvM+5iJn5SZwEvJDDwXjTMFfIx/vY67ybJ+nRh99ld1ZXinPfecZhpYNE6hjkhcBUuIkRn+RWuRb3zIB5jZlm1PooPKqvCVol3NaEFfwMd/nqbf2o+pr7WM0wg/vAziEeOpTPqn875f3d0WjR+bV55b2vo6f+QF0k+/GE4L3VVc9+zzq5u+vpm6jtzyL979v56FkedtImenlpnz/zfdaYHxNG1bfb4vrynO0PfTM/Pqs8lfzap+kZTJ/WI6VVj49+Gm+tCodzvxNpofz8kTsZjszPcvrp3cEt7Jja+sbU0+87/v8q0AlkBOy3rXnVgJ3QQK82dvUSqCVQCuBVgKtBFoJtBL4iyqBxhITbIkkdLIbwb/xMulvbW5tYCzs8j3ewWAawVMqPsw1sPmez7+oC0ZQ1w/2/Y96QIA9gCt3ooy/1nO9g0eJO7jFDnCNMSpQoefY1tYGz1jWBS0Rpl3/nI+RHH/lh/bugHs9aigjsOMSKtA7vEe2y8T8yXL4+Em8TsbxdEgwS+PO1KEd+RIws12TPO7By4i8YMx7nwGe5ZV6YTDRPLed4IcLkrvdbbD8Di+tAB3sF8bjKPbJLIDHCYzjo92JyeWdlfW+OEfaolWuQYIfVd71/s96hi6bjF548J3lPd/7/sN4i93X39q9DB9T7Eq5Q5ytEXYS7aytboS8RjqYtcghlrPBQmcHkMF+y5EgmZ49dF25aUTqMsLmaBjYlENOehwFOCZ0xriIagW9xlALmTbjH8YbBnYagNCnvdrr0A/oCYrRPCICfNGzz9hU5PM/HzSghSVM7i5p3LsKuJgbBi082054asFv8GGDJJf4dmLJVQIfgiZErOMJ+r28WBZv3Ywxtr9XX3qpvLa4Vm4uLuPRqNdj8j8BMGZMqYWFhTI9lQCZ4LFyyj4HwzQ2aAxsdBZ6LmfcUt7IB0VFpaFHh23LHTWt7yMnjnIFUpNl6KCbnMK7BtBgVE8v+q5H4D//nd8te3gBbgN6PP/8d8rJU6fKo488hpfYpN6CsYROL7iQbQjS8XQJp54pCd7oGei4hTecaAfPoj26EWPjnGvGUXbMG975zzyBDpcV8rTpcwO20IY71/aoH54sgFduoGF9atE33geAhmha1OUHe0vAL96k4ckE43oj6SE0YG51jSM2Mlmef/VauXpisixMzZdNxmWSMTUE/Qg7XzrUA87ffuVWmTp6upw9dxF5AZzIN313GaCi0KsuxkIeqCuwoj4JMFug9hkNCiAp3gfy50sAfq1LSPSQLRm0kYCY4GM+Q6aCfQqfxH4ecfYloH5mn6HUvJ9sL95RskAV83fgUanGEXUk4TvVAjkWgoruBhrjwq6sgp7qka+tZ555Bi+yFQoC1NpBUo8yx44eDd3IsVQXbCseBx3f5b7nApxRFrjw7frHDGSR+qJ88BKEJ4cn5zXPgobvW8pmd4MXe+Bck2/brLKNoQ05pk5VfpITddKy3DlgNfFusP4oSJ5npEZ7OUbp8Zty8dmYS/EDvlOeSpEz9Gxnm/70/UMN54btOMMJZXxPBOwcv38c+5rUR8fY946A6gj6oKxyXIUKYZc+Ob9sR9nIfca7c2zUk5wzlWZ9d1jeJO+m1KOkkUyamzL3WfQfXrM8Os57KcaMqvQbJ9ORMjHNxhCzM4du3771jtXV9efwNP3a2fPncqcVB6XpvpTb1Ergbkkg3z53i3pLt5VAK4FWAq0EWgm0EmglcBclUD/SaxMaGBpMc/OzmhqbGMNrfJxv+CHOdYdzLDOs3lfVU0Mwy5hPelD44W6+H/XW8/CjXiNOjMoYQDRSZg4dCvDG3fi2+5uxnG8AYBYGAEaXZ2mYwgCDpsuOBhDZBGgwcHfpsczs9DmM7AmMPp+nV1QaEWl8aJC4lDDowIvJ57WM97WdKg84jueV9xrwP5f34LUi4AddAQlAj/nO6Nip3vjkMWQUrnZUDqr8GLL2bOnNSMoEyxiZf+KT/zaj0juDx9jFre3+SYCxzhrx0VY31vdccrW8SuyxjTX6LxDJ8r4dYkFhTgnUVLnE9S5L4wiq7nUcGOEaeZZxPD0ERkzKTTkps3rtfZVdFOLH8HOvfS7eUMtFHcQU5wZwqHVtyzq1TXXSct5Hea5NkdcY99q11tGQrcnn5sm/qY67wKxyOHz4cFk4ejwAYctNTc6UmdnZMomhabL/zoWjh+eirVpfujXty4AMr/d55l6jv7YtffXJpYjqsbRN0qp0I4Mflq1t2J9r114uzz7zxzzQQC/l5s2bZQWwbOYQ8xQ6QbehJ62qt9KrPEVcLIAGgQvpV1kKANRy5nsM78wpH8OHZet9bSf5l7f01rTP8mW+yaW6Ae7YVLgt8Y5g7ujdyW65wa+vBXlyirpcbw8wfHLuaATff/rqtbKyxU61W8xl5rleYwPq7rIxx3WAzauvLZZ73/kYNBPESn7sJ+01uiPPAh2C8D5XX8xrkB7ZDACsxv+qYyDwJVA8xtmYbRNcx7JTiFc5ROXmh7SDLveVDx8FCIZMXFoZ7xNeanqjWqaOYYJQochBrdKvdLwPj1iUoLaB+1B4hn7jG9+wFWSYHr+CZI7D6dMn2SRAD8LqBXowJxLQq6BL6rtt1fef/KmvdZw9mxzVKMe958qL16Z677keyvONzyKDH/nkoF7NH6Zd60onvSFrW9Qnr/JW24s/sFBEcCyXhsrzAd+1DbXCFOOtUpCk4X2dGzVvn3ZTxnyTfL6RV++DBnQqvVqu8uq9yeemSqPe13Mtb5maN0QLp8r4vUtIhM725Mx0j2W1V5ZWlq+wOcuU7zgYkbgdraKWVJtaCdwVCbQeZHdFrC3RVgKtBFoJtBJoJdBK4K2QgAYQn9wcafhEm3gyPPfcc+XCvQ9s7exur/PR7TLLaWwh/oCeH/R8sO+xfSLWjzU0HHul39kqU+MTeG6k4afniIZJmLMaxaT40OdjfZRg9ofmDwN8dSJ2jnGyJvGWKWONwYUhOqqXE3FzsAgwVNIA6hP8fwtGNvB42sL74/i5C2X2yPGyjnGdS5c4h9FhfzDuWMqWRqdBsfUiwYDnPMJf2zU0NC4TWMFMsi/wqbHKvl/x3N4Gz41nTcTqkW5jdAsmjUz0ZvBoO8oSvfn1lWXcGGxbO6T6VXA5LF9v/4wpnAD2iD1GB7rzR8bvu/LQWZYEPoQ3xXl2BR1ZB2xc31jf3dra7KxtrGPIJhCDqRbg5STjo1dI6WgCMz7I09Q3/hjj3gckc0y37Rf3Lq805pF2sbpiXKxAaIb4r0aeWcrUew1LvS+6GOmCosqQJ3iu5ThFI+Y0Xia2Wevr3UR10gFIOgJgKlAx3FYtX8/1mSALNWOsOwyufIdHDWPWFYDB28tlp3ojnr9wqZw+e67MHT5a1vH0GhkHSCX+Xm9ljCWVPSQ0EiDaIYCo8XG97gQL0EcUQ+PXdoB39nVFjyOnVALECZaNog+diYyZtYceqTOhHei2MtKrBVaCFtHrIjl3wrhWEIzD7/3u75Tl2zdpVPBruxyamSrz8/MBgBiHSiAk+k3Z9PhKOzh0PISpPABO9AQE3HX3xAHeXrZhSm87nsGPxdOebpjxeeTHoERfg1uBE58xtmMAY9KyPZPlneO4euaYAc6E3lDOsR8hoHiXWGrOzRRYtrWLfIIEvAqETx06WnbnjpdXbn2z/KvvvFTmpy8Vl5ZOTPG+oermoFOefu6V2MH2/nc8AgYHH3oJ0b/w6pEsLCUoBr/wJW/7vDLfQ2+Qa9VdRjeuwwvNVxwM2SuGJAA254keZAku2VeUukmQ5t6bBlSiojoC1kw+wCj9FQgMryvz0eu6HNxa8hWersrFPxKEpqgLzJugo8TRJ9qo8eJcRvnii09zvMj7dsDOmQBhyJ5ldshqolw8f4F3G/yqhwApzsWu4CLn+gcOZeAhb74n9ygvHx7x/pO30O30flQYOdbRWWhnv2OJOXTSeyx1S6DKI+DJ5vdHtEX7+MBFf6JI6G7+nggZ02l+xzCWEI9fAwiz0THfBbYhaKlsfM/tj6kU6YfyDpnRTl0myqNIztGQLv3wbKv2J+nm/HbMTb7Fg1/fVdx7OMYxR5370Xd+kOTBFPQtRAr94feNMTD1qmZJfvyRSA/dDv0z6bEX5Zr505ziWf0hDzm3k673gs7Bj+/HTnev2x3s+h7wODQ7P48nLFjZLA2k3lRa7bmVwN2UQDPz72YTLe1WAq0EWgm0Emgl0EqglcDdlEAa+LWFUYzMr3/9a2WwBeIysreMsbLKM7+wwT3IaT78NZwSYEsjYGJ8qnQnxgt/wS5jGL/EQEnDAgNEUEAwxu90oRm9EroYcIJRLmfbwZAOjxMKUCtAnDBKuMemSM8zjTUMmg0s480BO8QRo+jQ0RNlwyVBepVAU56SLw1P44SxGIs8DZcAEbBmDFatAaFBEgYNNopnjRrrDhsqysR7k/VrnTD2MEoGLPHEe2uCanMzMzOz0LAQ9uPd+ETsjCFvEEjAhtHxvc9/4d+d2B7sPApPT6yub57e2NosLKu0z6PIYsT+uwlpsA+wI7jz/7D35rG+JNd9X999efft782bfSNnhsNF5AwpyhQXSd4SL7LsWEECBAgCGAaSIJsDJ3HsOIYdB1CCwDEsOVCQ2IH9R6LEhhMDkiXZohJLoqyNtCTDsjzD4TIzJGd9+7v7ks/ne/rc+5uRLJPmUBSNrvf6dnfVqVPnnKru2+d7T1UZSbYDGGZEnRFm6lsL9ddi/doccC39FSBntI32Un/LYyvObWdtY1umHhteW8cUR3Z0qI/tp43GIzT6evR8l9vGbB/N0nYbfbasrgtUqjarby0THLM84wuXeZcdPne2tjMN8IEHHhzWcSCNrqnF7N15UGBhfVhhofjTRJNdOn9uWF9dK9kcnfDqFJ4z953vw9IyuwB8X1u37VZRiAVMVF+dgBHSNa11P/0M0WM8Q1rp9PnLyLoWwFOZTW2r3Iw/rG/dTi2DIK/rN83W8Vr7B8SibDbJxzR7br7mHeePPBeW54eXX301IGSNC/QHyGDgBMASHJsHmPa5NuKseTmVNO0IjqGrcMS+wPoqawsunx5+9XNMtXz11nD7YIFjkcmyK8OdYXV49sVXhkff8Y7hIlMJta1jp3iOYDs20Ayd77mvjfAzktBphyIdgmqCJEsjD+3iUa+/6lPrdrK9Tm0Lz93Hfa0dMlZAW9TNKNoCxqp21XVslZ3LbvU+Evi33NS28myeZ6eoP/eZZzO90nr9nvK5c/OJM2c3Mq3XKCNTy2/d5iMvZWp9fG/Kq+/72nvrd9vyk8dsav5d1uOsdej8Op/oVfKoE/2AzZtv5Y/vBtoyeiz9NtPuLG3L5tmoPX9HKbdH8ka7tczWbZlbxuYnjWCk5QJlJsvezMf7bqNpmmffW6/t2Hmz7TVfyzp/9tzXXS79yUisOj5PbspwhuhsbHiGsXYfINzZ/HLjDUKdelGjhnymNFnga2GBKYLsa2HViedkgckCkwUmC0wWmCzwm2SBcvDGj29dAS6Phu//S//j8KvP/NO97/v+/+UWf/G+Bbjigv14tsQiEJaDD6NnI+zCx7xOE04Laysts2bQ3DwLuxOptLvttD7/hj8CTzqhJD/sjdxaXV/LYvJMC8wUt9OnloclgJS9OSJbiFyKMzEHqIaT7ALqOtR32MnO+Jv59dPD5XsfZS0iolAoOCI0qaIxjHo4WW+oopF0gm3XiCYiTGi7pEJ2nCblMZLFNW3UZbRFyYm83mcqGHwFvqTH2eTSKIzohkUO1y9ePO+8vHj50iDu6IScONHqb2rvRNt8eUlXSAOKUs0P73zqQ8Pb3v7OC3NzSx84ONh9P87tWQFJHUv6h9PC0SpgJTEWAcRsx50G9wAii6Yi5fYOiRgjqYd2K3AM+5PnWk461Q0cNRiqI0hTb0jpUzI9tyPqOYTYTxsaxbNDlEjsGQtIfwJMytAyeiDthy6RIjqwNmi7BVj0TpqCG7qJYymRGO0E69RqLft0LlEbWY+L/t0hyk6Q4t577x8uXr4yrDAOY1pcR6Ox5gFyXWB/Y+PMsIENzwCSdTrWE4Nqr4rAKf2UN+NM4hGQlF5HWXsuEPHoY2OedQUhFoy8YlxmJ0fs5WJ/mJ2DGujsc+B0yldeJnoMEO/hxx4b3ve+9wFArwPcXQqIZ5Rfng+ekTkiUUzqboJ1kjatpKz0CzYREos8EBtRVoQln/km+1D5tWGd1dk+lo8UPg/QcchxEfCLouHjH//4cMT6YzzQkAB4rJ0qfdDXKCf1dRyGT/T0mogi1iOzD+Wxi5w+k4fovbRxbthlab+f/kfPDutnLwwPPnBPplj+4rPPDzcByz76kY8Na0bSMUYCaDgqIrf3MEOMjKeMo7KL5bwA6Gvsx7jU5tZ1vSvI0YubjDn1L1ANyaK/5aZEpDpm3ZzEfoWf7Zgy/qnnre+bA0ExozdJ2rPo6pxxRF3rlJzWo6Lmg6/XTlPds4/RQdnmed8ibDaUeAYA1V2DV3hefWaXQjM33H///QDApyIbTeZs+0bSydsoJvuaZhN1VaAd94wjZaG3JUeIirRrWdTV5Ln0qHeC6+xZpAXN73I3MQj9yM+y2D+ZtEW+etWTTHMjne3JQ3zVFBhXvtGv26fAELSxjnQ0Hvn93fCGtSfRl0KeC9qyv6kjBmu0bK8jZnXb9MhApC3rqFOeS01HVultmS2PAuZOflUeMM/SjMWK3Ix2yKeM1kyE3FivbdZ2iwyUdT4LHMC77JrhWRzSn9A61ZKm5gHJNoZrV6+eXVpeeQLbvJ1mmH+7sD1GOyp0KTW2O50mC7yVFpgAsrfSmhOvyQKTBSYLTBaYLDBZ4OttAWYn4cThNXzy539ub2976zp/gb6OI7EPqLWyy7QsnAQ+0esj3elm8eVxbHWudDpcGHoXIGtlbTXgjBFLrg3Eavaj04IjDPC1TDlYzrC9tZu6ezjUe0vyB6jAkXb9bB3+PaK0jgCjNgVwmAY3EM3jtMq9eRbpNnoMB0bwQ9ChQRyNqKMgsKKToaPifRwO7olbgWcBY+18ODWzF3e2fufryBvFYdIhBkSZ29/anXPXPnkCtiyyOPmZe+6579y3fOgjyz/7Ex/H4Qs9mujqf7XJCXikOedFLt6+95Enhn/nj/x7y9jk6TtbO9+Mr/eIirI4/D6Loxvht7DMStsrq4vD9vYmdmGaKXa0H4AlEjEmMBW9AIO0iX0naOS0uwAoNKejbZl2CK1u/lFH/JSDO2uvAALUk75T2xA26R/tZTKyrdOxowfRcR9ROHstAOOosz9n+dvn2dVuBByUoUAGKpAiNzTALKkn/U0W6Hec3H3vfTmWWb+u0yEOteNfHutrK8PFcxcCvBR4wvih/7PbKuNfAEsc7FhHmLRstms61PlGLwFYzx7yVremNZJMsxQgU/TSxPYgNp/5zGeGa9dfHzaIBvrAB79lePvbHh8u3XVlrC+f0rX5ee42lCFtolNfe+72u440s+UtZ+dL5zF7bxu2ra4eAs8L2PLFF14ffu5nP4UxVIpnkE0EBL52eRSSRQRkosVAPU7eI/V82T+2Ue0AjDN2WVAJsO0U7wl4M830Z/7xp4dTVx5gSuzB8Csszn/3255gGuEjzM52LBAp6liBB5hHpvi2LZtvxhVyty52peCt946vcYhiDt4T5Ef3sb9GM4VWviiZcm0Xe8jMa9rWNo7zAPehq/FhvnrLt4BGo7dK/7Zzn31Oq52q67XyG+VmEmx85plnhpe++CLvTQBtomMt99l1o4T7H7o/19GZ8raBz3u34dn2D+gf+e/wvjVFn1H/rictPQ6fovXelPw2TnLq2Sublg29lq5lkQz2VKbDyGf0cMO4lyVZ3ab0EOTe3y9YNe2HHyXNz3vpknLd9vedUPIKRLbM4Q83STN+fZ65SXvHbMjjnyKmvVFf5Q0f6KpdVeBmtt7ISwDOJN/YFDrPpnCPrLmttusyfOUtbddNHemr+khZJ2iNGvaUHXevXLlyhp2LHzuzsfrYR377737+p378R7f5RYyMBzV43lB7upks8NZZYBpgb50tJ06TBSYLTBaYLDBZYLLA19cCft7XVz4REXdu3WSl9rmbuGM3+UA3gowP83zch64xDj/IjU4SMEj0As7Z6trysKCzRnTGEtPAMYpJIAAAIABJREFUnGKlA+13vVEJBIkMi+w6ucTW9PhqAdTu3Nkabt28ncOoMo+tLaYDAtyw6DzrYtG2dU6fH5bPXCAKjWiVMYpLp1PwSiAjYAZqOI1M38pDR7fiQk4M3I5ScnRYOMzTITEixEPH0QXV1dHDaCqmMAlCZQpj8ln8BQDq3OLy2vnv+/6/sv5v/Nt/ZMaB8VPx5HNRF84jBkzD/7wfqYtXAxp4tHDw4OPvGf7L//rPAzAsf4Spqb+HyLEnt3Z22eRxIbY3auz0uVMsMr+K3ReziPuZc2cBe9ZYm4hdPtGlgLB9wLPtRDF5du0x9TWqaW+cgunUSx0zp9zqu5Yfi6OK8O2wqf9sajuVAd7oxVnHwxReVqWPvDa/63rWDfZo/ukrQFYoy4GWCehUT8vzVoDAJK2RZTqm4QPvOKSM3V0Aw6uvvU6/HgRkOn/uIv3JAuZApq5PZgSR+jkN0alKG6dXM5ZbPm3HKInM2XUQGQQLjMwQs2i6RCKpgzKMeuc86qWMHsrVZx4Mrsshbr3d3fWTn/z54erVq8OTTz45PPLII8Mjb3t0uB9w79IFphQii8+VEW8e1pNf97PlRjV1KmCUqDUAY8EJzyqs6QIOQe9aVbEXlcyvabrS0BYIl7rJX5rWbYlncWmR9e2Y6vxDP/zxYfs2kYncz6+uDwtMV3XRfftaB72nH7eOiFvJ8vFGHUy68nMAbIdLp4YbrDdmtNg/fv6V4Zkv3Bg+//rO8JlXrg/vfPqD2aVxGTtXwFqBiw3cGWHX1wLyHbWoPC1/pp1iC8G1BfT0AGtDHsBV7cN48VB31zAUdLbPD1jPLgcm9p3mO9E/DuxiH9cb2+Wd5e63+6yZCPaMzbQdfUK+h/1t9N+JLUpvzeWhPapPGRd0mO0vRYeS/fVXX8t0+NusqedYM2LS51h9AUiGuy/fFdDMacNO9fV5cL05+zJt0rZRpZnm7ruBsh6PbiRwPD4ZnBV15ju8xq39Y6q+0liCk/2erfsQjD9sr4A9dayj+1l5/d1yXBtaNIalzxry8nBJo461QH+MEx2ih0g1h1MqMXds799S/N3i2NPuyqc+0tvvyYEfFDz/Pvvatw7/eGLUn+3aD9K3rNYIDx8O7OiRyMGRTtb9+y7rjklH8t06y8O8N9/nGfE5wBYe9pXnfh5rV9V6R6S+ImgrDsEx+GExxirj4PSZMyuMgXvXN87c9xe+7/tO/Sd/4k9SRVrfVFxMabLA18gCUwTZ18iwE9vJApMFJgtMFpgsMFng62IBvsxNOEcusDUM18Yj20D6Qc/BGs5+xZcz7l/n+erm254Pdx06KghcGDG2soZjA6iwaxQY99L5se9UoYWsRcRudHtbKd/aJMLJKWc4mdt7mwA8a2BCRDfgdM0BjB0ShbJ8CnCMw5igBRzfOBBcm3QSFgALdP50pmynHaH4Y6GCTt9DJy+6VD0dflNk5NwOpPd9yH/2mntmkRFYd7C8tM46Lzhil9fWT5//yEe/Y/g//9pfgQctWOErTzGhYnAQ4rWwTeTYcPauB4Y/8V/92bM7+3Mf3t3f/a6DuflvY5m4KzpzOzjl6LqIE4aPeDisrBqlsx55XZPITRSyNhGOYAAx+kOdtV/OtOT1oevE4fjHlgurAEVMewXwbCfRfAGBBYCQXMPDcx+zqiYPFdopbds1jeWzZd6bPNtvnq3jdYZbSuPpVlnuxz5LNiAVLJzmBcHYV1zSA/KxLTcoEGxyvTynVy4D0CaqBF7awTYFwZyidoqpl2sueE6ZkTktzxxOtAv9J7rH7lXssQ1vbcsy5V4kDHKPAS34FlsDOsinRNSpRT/iAyMfbR5FBviTH4CWNePcndC10D704Q8Pb3v0sSzOvwwgZXLTChf6Th+l3bKh/EzqbOp7r23baYzKoYzRm3xp60mSSjr7p54L7+UROXl2rdd957OW9kEvbt/ZHv7fn/gpXgBMd1w5xTNbu8sKdMxR7iEohHkCKOVilDVtwjfnMhCXIBhzLPbPu2BYOzMcsiPrbVCzn/snnxuW1k8NO6xB9shjTyDP4rDC8kpIFbkF+YQBlFfwyznhLW/zTz/YeZQJjHFBXWyAcE4upHbyynY1xutaW0kPhYOL5JgxqYqHUxc1nbp6+I5UpVxTZvId1NGazdd85bLp2F9m3DsFtuWXFmnS5iuvvDR8/rOfgYY1HdmAQbC0N2144IH7AvK6ll7zTV34Od1THWYjyYyIFSiL/KNeXU8z1VRA5MHKvh9b5shLbvPus3X7WpX6vq5GPblJ/djH8Y/9eYit18+85d77zDnWfBeRk3qW1VF8ys7YGxsLWtkH6jjbdtob2613i7ChCvJzfABsz9Q277M2YBTzUi79j9sPP/U9eR/KO6DeOKajAzaXV6eWpe+73b73LB917npN4/gZzRpyeKEAbz+U8PJoaW6Vx+0KRrjnzp3NU+94xzvlxnHyTKfi9GOywFtsgQkge4sNOrGbLDBZYLLAZIHJApMFvm4WKK8A1y0f0kcH4D+7V1lX6Or84ZGIShwVCplZ51/dcWK8iXOBA8N0R32BMMFhc92ZfLPjTPlH670dMDYdoUR9wU4HjS//bcAaFpnHwXN5rd1EaR0ZbrEHyAB4ML++geN3alg5fWFYYle7ORbtXlhez2d+QDKcmSUcAtOK0U60lzWRIkzlx5kYnYw4GHgOCuq1AMGs86HMRkLohmW9F2hKD/UrUMGpXAifRP151mlbX11avUCExCXuN6h6G/ajJ3TiEI0Gplj+o61ypRHLdMfnOdBCAtUIBzi6+8HHhz/5Z/7bu4BD/sD27vZ34QW/jzXe7qJHmIuaCAZ8dWJMEFBTxNFUfmywwHpwq4CROmtOJ7x2TcyTdbmIEOuIkVrMugGQAhm0SQUbABgY8QIYc4SznQYiJICE/Y0jqh07XzUcGcmDzrV9nOLpPf+T4n8j6LHDiw6hZ5y0rSXUSkaGxVrU1UhGh9HDcdi9avrIK63tCQDgBwqSaH15Y5ThxrWrw43rV4cHH3l0uHjpLngBpDIG5WM9+a8QiYXA2fExMsFTAMjoHMeKeTXVi3qjs+uGrqFVRugL+NAK41jyeQC80DY11grgWICvPNXMMSzwoNZG7zChdvjMc89ld8LH3/mu4an3f2C4cPEycjIskGGFsXhwuBXgsx3xRLJQr+WWt3o5/j03IFN9pWXKXgILjm0BMSWwnjSCAUkYUp7NF6tXu5wTfYNMq0SK/cgP/tjwhRdeHIZz9w6H2HHt9JlBZP0QoLvsQjvYyr6BPefRWUff9LYIpykdF6kTObXEmoOuO3iwuRWw4MXXbg8b55eGC5fvHe6958Fhl00XlkC5VgXIlXnsA0FhbS6wkf4VaTAxLtTXtah8xom9SdSYyts/DXw5ziS2n9W9k3bO7qOxqWtLSUdLPCemTNe2KeRI5BVtJco2WTU+CzgbnzUrzSZBWHlS376ITLbPoR3VxejCT/3Cz2fKcDaWYLMJ833G2TBkeOihh7LmonW1Q4FG6mc/OnZlJ5DEq9bp7XZKmvBpiPD5Q0f01k6j6eDAf2TgHQmkFqmVycO26lo7lM3NyyYI5phNwqJ5L/SYEuS3VXed5aEsIs5eGREs8OQfXVxn0Z0rlTvrk1Fe8lFGVdfosq9jL9TJmQLB5pIrIWPhX2WjnthNkJG/yHBGDnjJ1zoynvd9b1v88wk5LjPPculmko+xh+8uoxEdA/ZjZLUOh7w9z/JKPfJdXiD5EERO2Nu3Xkcmnw+SkYx5VrQonRrAfeHoIH8M4eUG+H8X67XdA1J9OpHV8GANBYW16SlNFviaWGACyL4mZp2YThaYLDBZYLLAZIHJAl8nC4wfzvGe9vjQvorzffVwZ2/Xj/M45y5Wg2eZD3ydCElxcPhCzwe8GQEQ+NDXCc3HuhExC3rFOgqsMwatU9s2t3HwmdJ37dYmQSJEPIFN7PLtv0DZPKDOKaZSrgKMrZw9N6xwvcTiwyA+BY5hoFq3RrbKRkU9jDelkrvAjXY2+EN7nNg3OC3I1EnnRH7qGIeEAut6oM/cFuVZV4qzeRhgBefkwtzK0j3La+sXkYyoLxYIOvFD/nlOiY3r9XgYNaaxOBbWLt7z0Maf/nPfc+Vwfvljm1s7382mBR/e3NpaduonEiJq9YVyCLDsM2WqI56MjsKNClvXJAIWyw5niX5SH4AgwZU9okcIeIv91Nu8RXYZLWDIFduIThGvQ98j7UyKLQCY2j7JHH+YJ48DImusYypbFoFtJOomjjF50KT/qjh1Wo60qWiOp/i3jrVyGOmdsUaVIyX96ly2AhZ0lgX5nF7mOLzJVDTXYrv3vvuykYRRjOqIwTMFyml0y0TiEI8EqMhnPjbyfjlO+ahHxK1rZdQOZfs3ggTKHZkDLgCAaY8RELLMZ2M2yVF6EywDKnzmuc+xO+HW8P6nv3k4y3po7l5pEtwse56AEnZLTeMr8CCEMz+UkRbGemlNs48yMm68kWIc85GlsqJfCsd7wQrLE0/DIvqCGq4F98M/+nE6hnsi3Jwa6bpjh4BWAgvpNPWzHuM09hE0hCaArvmOQe0iek5fGs14QKSooPr8GgDZOVqEZIGxuc974NLle4iuOwutC9TzNpA9egigCA7nDN/oEgVKP4cN/4PF+C7IjVJSV9rYShCCMnkw6AOMCJyIgXWkkv3p02W94EujDYX2/N8RePKTxlRgm61Xmm3TtuudVDzDnzY0i8n3rOIaaSjQ/SyL8wvOOA0671mv0fvSlbsyxdKNUwpgKt1aBmVVRqd3OoVdQLbGJjbzH/k9fblt13L2uaLsRrlG3aSt59j+q2Re1zGH29i4ZTkpx/a+Wvj9YZ5AeHUMABvjzWSxtnSqphYMnQxnkn0jUKQ+PeaVyXunZzJ6Qt1TNeXRbfoMjaqEt4SW+66Sh7/XWu4wmflROlaGtMpctjjpS+VpmaVPf3L2DWt+A+72gSk0CkRZ6VLytAz2uX1nXdsLPWgc8h5iI/6Os7Sxv7dzz9rK+qWLTCf3XbebhTxLzunnZIGvhQUmgOxrYdWJ52SByQKTBSYLTBaYLPD1sIBf5aNXoiviclQ7NzZOnbnBhzcBBoAoOIoQhM4P82UcV5N/4fev+zpWfrTrjJRDgTNiPk7PIs6JDpmujRFL2wAV2zj6SzjDL1+/wZSpjeG+c3cPK+cvDmcv3z2cOs90yg12EDQS5cy5ON2gHTgKo5jIonfqGkE6gbgY3BZQdoSD5HpDTgfU6QLCQAYE1cGkzKlUctHl2nfNHutLaI6OEJeRc/S9KgIBBxwnRJxBZ8Xd0XRM5MSxTIvndvcO7ob7JeR8hWwAsvCEi27t2GQujh1I8uMJ2rI0iDJfWAVTyx54+7sf/tN//ns+Bt8Pbe/tPYU2j7Aw/7ICameBBRMOFaJgV50t881WNu2gM0nztqKDtEQU2BpRZUaEiSc65ZLlynACdVBr18tF1yziWGH3wTkBENuAd0A09aaNBRZbN89UkU+eddJoHGzPaVza9ISGHqLMqAojcGJLJFdpVY+TR5+V/e0PSug0I44cdfavkRjm4w6Gr1Ex0ncbntNv5McZde5c6qg7UwBv3xxOnd4Y7rr7nmGZSMREpdC248WkTEv07dES01SZVmkycqzbEIywjZpiZin86WKGU9rJWIgM2kLZdXWRCfZ2qrsyFoBT7SmjbUZXualz0iHA2Pbwi7/4iwE6nnrqqYBjcYgFHZVD/om6rDGoniZlNWKnZTZPu8fBpi89d4SUeiSfZtWWx/b4Xj2drhqbypu+8KSMZYPqMwzEcmOnh2c/9/rwK7/yLJtoAFgZacjhrpxG3BjpaT9mwwhkQbgSV/DQR4TxmXcIxhSEqGfcYUE+5Ps863OrZ4YFgl8c8+xAwdhcHs5dvJgFyVcYa3mGAUflY8o4pH9aVu3BDfKf6BDdbB+ediHUoXe00SjrD5ZNgRxUHzvWWIsN00ZheYnIshxeDabErujjWmNy9lAfd8y0MccKOeQjFv98BgIQ5h0HyGt+bE4+fW6kUI8PAdLPfvazw8svvzysr69mQX7pnXrreHr00UeHsxfOR5e0F7lLVt9byuYbSXDM+6xBpgGQyjbmeW4cG2/ua8ew/xAlOiTyC30c09Jq20R7aWuSWquzF9qaH/QTt+l069TYz/NNXrfJFZbRJsjDO8EoLPsvz475prQHXfq1ngFL0jfYLZGhdhrJ943TT1OH+oLTylUyl9xem5SBnyVv7n3bUNdsHuQaV1yTus7JddthlCtUyo0e6j+mHpMin0Yrq69972Y2KctohBhjKVVs96a65nlgQfqS0cT1+LsXVvx2po/n+d2JjBc57rpx48Y5fp+7Q4k93cKE/ch6Ok0WeEssMAFkb4kZJyaTBSYLTBaYLDBZYLLAbwEL9EdzeTf4FTh714m+uYpfsKXj5QLUSXpXfJTHGcHZ8CveL22dCx2kBpv6I946ggSZmYh/6If8FlMr7wDSrONIn7ny4PDkBz40PPDQI8MZALJD1obakydlAmRsg8eBK6ATQbvlOOM8GE7C575OUhwCPLdusxwlynF8vA7qRNs6NUZ/8T+0wAlIV85GOzxxxkal5Gd+dANB2GNdqJQvsGRyeBuJcbDADp9n2a3vyrlzrJ6ehZPmttQb6TQNKR5oXY4/qV/sdQFRbH5xdeeQaC7qn33gsXe967/5nr/4seu37vwr7JL5QXbSXHfRb9jZCdQ7WkKO8Ma9Qh/tXk3J9MDVqkmCHkZQ6QjDN7Y3mkwdPOzXzVu3U1ca+8Z8NyRw6pbXAmudCgQrm1imbW3XNmdTZIn5dRZPojC0vfVM/yxn0/IcetOk1qvP3ab3uQYACL2O8ShLl6mfxxED6tatWwETzpw7D4aDbowvIbXjvmHsLjFI5+ZqjS8XvjfN6iZfwdcAOohnWUkZ0mNbKM+JnFq+nObm5Xk0Qyq2vMVlGF597ZXhs597bnjf+943sENq+qKifGq8V0TMCBSmD2ocl3xt3wLAHLvmW8czoz3NKEPJM9oxuglNvLEvdamrr4pvwHJoBUoFVQmBGX7iEz8DTy5WmWHMmoEOVXGQeZ9dzu4EK2B7bGvre2AEAaDwQR6jGqtLcPopY3eQrKHHHhUAbwK2CMN4un17c3jggQcAhZhWyL8FFy/cx8bwzLTGsVdm7W10lW3aL6Z6X3FBG6b0JO+XLKBPG451aQ2aLT4FRDQPp4gLYgnAQD0+Y2gYe1lmO/VsWOdkmmVFemkPAcTx/9jGrx0nyiYQ4rMjyCio/Uu/9EsZEz6vq6urqes4P8tup4899phVkkrWkl9d1MM2D1jF3vEgoKfebafQU9MxbW87jltf7RV9sIe/AhqMtLxTX8vPvjUljzqC41F2zJultZ30AG3YT/5+qbZP6tdUxxlZR/5UrMT7yz++xK7o1v0cZULBGOS8QL9aNc3k2Sgdva++q/GgfNHDc2qOY3bUt202tg6/soP1Wh/LlEOwtfWdPcujWmsuRS+NR8rH8SnPbtMzUiMVtbGtz4R5qcfPsYr3ZxgX97569fW72M3lDs9aoa8nzU1XkwXeUgtMANlbas6J2WSByQKTBSYLTBaYLPCbawGdknIWZ9r1K59j/mB7e/c20ypvLCwsbR6ymL4f4XFgIXDKmFFk7vzFl3mqCxwY/eGHe3IAbZw2cohTx9onTFdjzSXID5gGuLZxbvgj/8EfG9715DuG++97AGBmObtW7jAzcQ9H5xBwRBDDKAUd1EPqBCDAcdIpTBCCoI/8FNhoIbxyHQYdEs/x5yjfx+kuZ1apyNCxQB6TgFsAPdoRGnDqTTk3FI4Oh2cdb53UOG2gfdwWD9gFQDgcThHdcuH0Bh7qIooC/tGyPLTnGxNtyXMsWoACE6/tPPr4e4dv+x2/a+Pipbv/1ac/+C3fefXa9aex4INMqxzBMR3lRTYHXTyiHzQtjhCgB9yVS/t4BqyTfZIO0wE7qJm/aMQGoJCOtE79OutGmWJXIvqOdnTAC0SRfgU1pDU5VVHHOjaK8VXB9ko96Qukg5ZFdNqRs32qpf2OyJFfojpSh54a7WzP6ESnh8Y8x2eipciUVxxD6plGnBb97U8datZaYqx029LYvFGGLvItQHYvY63t5DhyepoRQtYXCHT6llFKjoNVbLXMRgXuQKcdAqYKoGh4bYBepX0548rnvfJ2tJt8TQLEKma/lB7qCrDH4ULyxUcbQscz8PnPMr2SnVyffv/7mQ5aC63LS908ql9Kb8ef9rRc3ktOaxzpui3vtUXyEbzytafSvTElUjBZ45OsXupEO47ZTH1knCyvFHi6uXU0/Pw//OVhOHV2WDh1hlAmNtjAli6jZ5SboE7soADkMQ8YW2D3UQ6UOZbXceQT42vFNl0XqmSWF4DZ5i3q8zxv3Rre8/hjw6kVdpc9hCdtZKyoZ2TXHsXDtcZ8zamqbUZngREJSHUq24nhcXUM5il3j23XuDIyMvd56B3nMghXGoM/bTmCDw9HnVFk1naKEgGpmD4Znx9trrXdHVWmtit45Ts24vsu9VnnGX7++c8NL33xC8g48AxvhM42HBMPPvjgcNdddzHe1EftZFdgmA0X3+LttYdTEj3XtFTk4PnNOxYGsT315c9alNxDr+3C+biB3Esze/iYSj9GHo9lZTOfH9hUnn1OG/Uu0aBjfhRAZprxvRB7cW6g06fGyKs8b6Me6iJdKsEndbBx8qDPc+PDSJsN+GXMUafex+ZrOxod5UvEJcIasRpFHZxvkDG3/CjZHUEe7GYTUNP3XrcvRdUuckcLlGN7RWfbkZtz5IDUdJwHvZHBAoFNm/5DRv5lV2N1sox3/NLRwd5l1qW7gu5fZEg1QNZitNDVyPRzssBXaYEJIPsqDThVnywwWWCywGSByQKTBb7eFvA7uRzFURK9Ho7kHeEo3eZDe6vWoMLpo9AaWQMLRwG3gXugA5xXUz7YcVpMIjiCCwJkfrAX+EJEyOrK8OCjDw9PvsudtYbhVrCkg2EHEMwFr50OwwoqfOoLeABe4AhaNw4CbdkG/2lbP4d7paCeme7Q1w6H7R/gTCuh1DpPOj/taAS0GN2DTIOBl2Vd3ud2NuThDocCKUaDMIVFW6Vt9GSN8PmzV65cOf3R3/G7F37yR3/QAmXTDxxbkZqkA3eckOJofu9g73D4fd/1h4ff8/v/0DdfvXHzu67euP1dLBezrttMxI4WIsKMiaoHrOZG20bxCAi5ILhJmyin9jYr9kgJzVFbZ/CQpjxLa4SYQJDRZFs722VH8i3TibRcfjrKOuiuCTTLU9aztvLeupXKhtavOpWvk9sjrcusc1KveHSefS8d2tBW8bBN86pt8snWcTeZZ3vHNI4L+l+wYPP2ndQ7fe5sACfWisPRrmmi0htlB/bg6IInejOejaBrvtL4VIjczI6hEPCj5CzHtvNaD0G3TtpW4CNlYVgl4e8lfWKU4q/+6q8OF5lCeO+9LHiPTsX/xOb2y97edvg4HuQrT8/y8tpkW22vlqesleL8kL9lqtjJe8FGgQyBGXk63o4jCL2mLR6p4fNffIkpli8Oc+tnAMYYV9gSwoCq3R/hqx3SV9iQemOXpqiaLvtRk/ZsX7CoZBNsC+BMJ9X7ZBgevP9K7GW/uUB+aWzTctMWNU56187SofrC60S5aSfaoKXUd+MKr2r6IOOHMbTP4yf9Ud53Po9UQT7tVVFiVCFVvlfaq55H88q+9EsLKAkJqhpvMiL5PsourDOvi37vWe7z4OL8zz377LAJeCrAjZZ5Vh0Pjtcnn3yyduUc+822+Y88vv+MpBUQq8ixvEcshEvGF7bw3GOtx5BtJ/HuhBP/65mNPbkVWPMPCALHph5vPa7M67HX5bmPxc2pOvabveO7JuCX144j5UIfTipynGe+KWA0fRPpKN9l0wHbNslT8ypTPyPmc5vU7zV5RR8KPHdyBMClb3NOuyONtF1Xcdp+LZvn7kNHaNPKqMY5uccAXrXbdaWZlcV7U8vJVe5tU/Bu5A3umw1bQkdk5jIdc4VGrhDhvLK/M9xOpTcrNWZOp8kCX60FJoDsq7XgVH+ywGSByQKTBSYLTBb4OlqgnIg3C4BTkSkam1s3cbqyEd2uH/kmPs7xyYjJwRnwL/vxl/hOd2qgIIMJVyMOyiFRVNn9ECfDj/iU4TD4IQ/YY3xVrl1nZk8MiClti/Osf0UZHMvJQcQ5HHTXoZEufHB+dBKcRQiElva81xFWLqMK2kEKHfXjrFE/068iN0LrkCFXOdTw4tp7IxJ0PbSOGiVyQ6eQXB2qkZ4ZZvUpqKNbpHPri8vr63/hL/xPi//Zfzo3/H8//H9TokRvSiGPL6gQKOeUvqVVpqN94PkXX/hOpPqWnZ3dde1xuIuzuEQMBmFG5IHjqSDOHiDiHt6OSdtF7hHQAPmKbXS4zTeCp87Vh64HZ18tM5VVwGN1dSv9oAOpnQTHljgWiKCy3yGNvY22MmlTHWKnxcWuo4atKU2Gn1iIzvMcSITRUkICNc0WqwhEaGd4wXF0XnVOy+7MHyWf/oTONZF66lw7mNbra8/2hWspFb9Rb9EJuUP78ssvxQbnXazaxe5xSo2KK8cbOUaQqaaB1XjVHpEBxQKIuCYSbTXgorC5H/V3hCTFEAAROul0grwdM0alaU9tod10amcBLfNY+G949ZWXh2eeeXb40Ic+nPXS7LvQw991ihaMYsMupTPPGPVK1mq+7ZL9NOi8RPEgt0lbIDX8tHvd54IfXc+zqSKW6rn1XhnsFoFFgyQXl4kIBbj6uz/+CaZL8/ycOU3kJ2M5fV31fJZMAdpy5gd9dSRwSZEvGkyTZ9bHSNMJSjhu3MhDeyEt+T5JBSweMcVwbW1xuOfy6WHNKZd7u5FNHNkRqq3VQSBTbgIQ82lHveElP0u0hRfaAhpBZ/N8o0hnSjn3nvvyWyUvAAAgAElEQVQ4zs+4sLpvskqxbnSGj2umUUkL+AzmQeJaADb50JUMCkE+feV6gf0+UgYjy3y+tcM+UWlffPGF4bOf/WzGkICYehrZuMLulffed/fwyCOPBHjraDM7rOoiDyrtA8Tv8V7eAUjX7lFTmyNnpjZGEkSlXo8DhAiPvHvQJu9E5EqkobpSbj+7UQMc846N/aEt+Uo/31sm3z22J221y3tdPtqKfohNfDYhESjLLyP7n/vQUdMybW1SDqOE9zjcXVS7pZ+RK+2jS/QZ6zvubMMxhuDHbUpb/a4eFPH+cO28XENvneYD49Bax2R+2Ml3zIse1rO9vO5DynXZxTx1QOOxTuleVOHKD3WssWgEY/SGZ54L3yO8QyITXFLDMDx/D2KLo9XYeYWp5Jehv8waZOyeAa/RbKkw/Zgs8BZboJ7yt5jpxG6ywGSByQKTBSYLTBaYLPB1twAf465nQ9rF+d7xI1xHkmvdoTgHRo84HTIOGOCEuyEawWTUink6GzruOvKejbxyTaJlIshcQFhHUWeUNbwC6ARw01GNg0PLo6OjEOWAlGPZjocfYtIa9WFeyyW9KWU4EJ57ClrouHfjAJ26dmwEL3Rsmrfn8OCHDqj36uCxguwr7HIoWmUdnRb0naedZdyPVf5ov/ytH/lo6uPsUloOTjKOf2hQkAYWu7f493/3v/nYhz78UcGx38eUnIcKnNJDm9+njUUAEf1S/MMTh029tLdJm3ut3V1DSTrLTcrstbfVVwWomW/fGIly5syZnE+dOgUwtpjIMsvkYx1pvVZXz22nNDD+6Pa8tVw6U9Pnhh/dl973tc66ySrSt8Us//X4mN/tNX/v6W54yqg44EoizMFwlTW9tI/rNalj65ZGGdeCDascntVV/m/uN9vxaJk8t56eO7VtCkytOl0v7WJE6560UzW7bz7z6eeG61evDt/0Td90ouOxg1326LatabQTu2iESbftTfOXtlPL633br/M8m5reszSeOy/4LH1kYAohjcMr124MP/aJT4jvsmMlwJfjBGBVwMmUqXEOPFIijRocyWPBM6sj73VsGzhEyuQJeM7KaN9qR/vz7rsuD6eZIbwg+C0wwrRNy2r9sdJNvn1Y1tdqKd8GCX1vCIAqJtpyVD1eK/Bz/Pu+m+GJEQSL7K/wzIurxrx6Fu8CZ3KPHN2+ZS1H53k2mW9Sh9bbcz/bRo194QtfYKrwzePxax+nDnTvete7ALd5n5CM9pOfMrY8jn/BMd+FJnUySaMM9rH8+tk4lmckbLmt47X0LXvrYpnXnd88+l7AqXUzr+VHmuM6x7Twb37Npyw0jgMLx35D4/RT/+5p+q7fZ3nPjuewGO3u9WySTlM1L+t67dHvwVl69WqdUhc6TVcbNczIPFOpeXZW8zd/NrUMKadg3rBJz8jY9vTeehypbL9yrGLbK7z3rkBbiytKqMGmNFnga2CB+jPa14DxxHKywGSByQKTBSYLTBaYLPCbb4HymOKE8Nf+F1/44vD2J57c48N6G6eJKLLDZda3IhiECDI8B/9yH3AIR1ZHx0WkDUvwy1vAo6N+FnDWnDKZCDAKdC533T1SZ5pveR1Qkx/7gnA6qIm4gJOf+ov1vR9HQAehIyyMktA5iNOgM4OzRPE47ZBrJfE+6xPpS5ED3UmEic6S7SIHdEae6djLT7rip07S+NmnnqxNxQ56uMbD5hYRXNBKb8IBnSM6YokAu9ULZ9l5k6S6VZrb2R+EnRAmMbe49PSHf8eVP/Td/9a33ryz9W3D/PLji1Ta3dtnfXImiQK6CSAa7YS6gIG7LOFE9Ac2UXfP21vbkcHYjs63bI9NFQ6MsBmTG7llwXHquE6Za1+x+BnKnWJa0i6gGLtb6ixjx/VVoqxIsQ1rEu1t7xvjhhzaR/8LR0zjktpeS9jI+tSq/FG+4Aexqw6nBhkdyaqMzNpaXqPdYX9oYB18HAu0Gn4BnLhy7Z1uU31tLbsfEpMYm9CWUAs/aA8OALfXr15Lnxodl7XFADmtq0MNs4C3S6Pznql05KmnNMrlucdXyVrjrPJLn4BxkDvu1UlZTOGAEQpHqd3mko8tir8jgb6gg3aH7eGn/8FPDg8+dO9w+fLleka0A7xKTyKKjkcUaxy55jbt+YwYayWN3eMY99kUbBFAs6uMfHNcJ4/8bltZTH3ftrUvQ48aNqkErjkogHIIz3kWzf+lf/LLw83bRCCevsSDylhit9A59HC8KrNjVvnsc1HwTCFEQN8HAltJoz6C1jbkyFLgtjNClGzwMYqReLHhPe96B6skGhHFuMTWB4zlCEnNtrsAm/JrEDfpKN2RCbs7ldvktToleswxah4/ciBHZKiOg009c74DEq0KX6eBSuNOqA2Iat8aFwV05RqVHKPVOdDTDuySl3XG4GWfaSfHj+NWPYj6IdprN6DWtdevsv7Y88l3F0/LM70UPnfdfSXTK9VReeqdqnxlD0GaTLHEJkZaeW1SNut4psuySYXvSWWz77oPciY/iZOWGu/SX5ZbTLX0a4AvmDR/R4/CzLGmnES+u2WQnWTzxwrGVuiRYZSn+VWjVvePFI5wEufaiMSnjgPe2t0/2Jwk9YLUsWHyJsC5z0lHsfEcUxQb+LaBR8YJ/NAo8idKC0PbUqesv4koZW+1rpS+hkf6JiBWjQ9LHUYFrHHj86DNItM4zmxxtEHJUePButUOsqGLz6XSWV+dTdU/NMBLCju6DtmhEYHIvMzt5VdeffnS4d6ei3pCHRsp9IngMpnSZIG3wALjE/oWcJpYTBaYLDBZYLLAZIHJApMFfqtYQEcHR/TjP/Z3h1vXb+8yJW+LNZm24wTxte3Hfz7Ikbev+y/3+4ARfsAbpaDjEkeG8y7ThNiNkcN1xvyo77/449hQ7pEPf3gLaDX/AiXKMbW887vdciiqvPP6LG3TN53Ogc6GThOYRBwSabrcs1Mtu57OM75rOTJKTZmH0XBLLJYveBPnGrn1K5nmRfzYIljTKmgBWuH7wLO8mOpfkDbmkbqm0tzS4RPv++Dp/+iP/Rcfwya/b/9w/l22j6ctcKPzYjhI1pTRvh7qJo3RIF4LbJlvOrFf9YFRNe54J600fa3Tbb2mF/AwcspjY/1UIslcm0wbRR50bL29b9u03Wzb69n+kc46TSvNm/OKtyPBNcCKXrqO/rL8RIaUhF/zlXfbw9K+9lybMCjTHps/3GFXyJcHFqpGt1PRs3lYT/1tx3omy2xb/i3/7LUSV/mJLazXtK2XZ3nplLYeTmn12mzL6rpcCtfBe/GFzzOF7rnhve99D1MYK5rHvpptv2VreS0rneu5nJXDNrod63Udrz1MfT1bb/ZaGkG20AlQGJ3EEN4EL/ihH/v7LMrPLoq0ExAXlj75qaP9ZoCYzlMe+Xf7IZ6Rx7IjgByEpYhngXeKU0t9R2RsIMN73vlkMIaasitQHi754TtDPeXTz4x1naroe+g42k7Egr5JU1zORpn2WI4sPsQ56jH2PZZy6hyvyTZjS4WoegW2lH1PABnLzUvfALYt8rwvqgjJep3UwXeokWO3bt0Ybty4MVx7/bWMV2kEe02+i9797ndnfFu/baGMOQKOVXTv7vgu0C7dlmOwnwH5qYplAn6dlNVUfec76ESHFPBOX+KFahXP0Y9rn23XTuu6jo5+HRbPep91fvGv567bpCXq1DiWj7zVy2S/2m/2aUccdt+rg3/Y6DGvCtUXCE+avU7GmBfdaaPtI12u87YvsM08U8nh4Cs9zNf+HcHXshzzSK1q28tuw2tpmu+b6S03yU/ejjuTdMd2qrHDfPyM/yPe++zPkt8T5x96+OGLjzz+DubU24/pSxUoJWQ0pckCb5EFpgiyt8iQE5vJApMFJgtMFpgsMFng628Bv5aPXSIcjr/6/d87PPvss/t/5a//wNYCC17pSO3tuxKKH+Z+ZBNrQzRZO2J+7Pux7lQqeRnp49o/Jv2JrAPEX/A7wiIf937nj43GKWjvDg6uAWMevocc8t+6rEHMvd5OOQwiU2HR9JS2U2T9JaJaTEZGLeBom1wvJ2vo5I4fAgACd/BUZOsZweS9Ah5knSHuKTOKYcX1dvBPnVaayDnkTj7eKhFea1tbW0xtyY5hEU3+YwgRHg0MFteGBx977/Cf/6k/9+Cd7d3fSdTNtxE5sYGzd0RkBLPVFhdcrF2bal/1OdxzAWqcc9YiMpkfAABfUZBOmXWIRP4Ewdxxz7S7UxFnEOVeOqcaApOljr0VOxEBpHOrw22UVfpSOyDu8gpRgPSrgIcL2BvpomNvYoG0yKlxIE9fqLRRGnCmXk0BrfIaI+pTETcSUon/YgTuOOk6TC6l0+vryFQ7uBseZEmRJS1RhwZ6RzcLlS2Opzxo58UXXxxeefm14ZsffjvTK08TCVdrkGmPJRo18i08mMUqvbIbWRcZxwaNeDEqx2fAB4AmkJVxlbYEbl0TrNbMOmKtsrRPXUemUXgtPz0V+fuHbQhOICl9tjt86pM/N1y4dH548j3vSv6OEVIsfA/GMcoImIg9EjFHPeu7rpTPBRIyzRFbaAO1IE857Sbbj804l4YQOd6lsaYRUBBGbvrbCCajfbynSG4pd2rl8vrasHb+7PCX//rfGZ594dVhbu000WQsbyT4Bw83jpAnEhc/7u1D/8mvIpSqfyMDlBQgJ+UCaoBGOaBXZvkcHNR6eyuMy1PnTg/vefKJRDg5BncFe9DFxfQF0LSPgJZjOuvALdA+5ah03FzZoOTxsZBWMTMO1BZdIusoe8YFPMzT9j5bx5s1ZKzChDXHrIomIz9uSNrFMaP+I0H40GQiB+k9+Clf0dvGHjoJjPIeye6rm5u3hy++8OI4JuUDJ9pV7ktX7hrewYYnjgH7W9BPHo4L3xe+nwpIpyWu+32trh6+CwXoEs1FPXVIQh6sknvraUD5qklO/kAUI1Etd3dTX21W8KdSOqbUUzkRN7YTRct6Z/InP78vfO6lyei1Jlzgn/6XwXjv82eSVlWN5Ov3YN6ToJ3hKS/bRkQj0/LmgJ9tmRgeyAeH0I3vL+gD5qED2akfbWfA0SCAFoaH+te1bZraptpDsDBn2lQXf7/Yril8NYjXo561F0vpZl7nN02I+SHAmMjF5gVtv4vzByl+FxAhebS8sMAQ4Xf23sHS0x/4ltN/42//4Km/8QM/MPx3f+ZPwYMgcJIsfCN0Ug/bndJkgX9RC0wA2b+o5aZ6kwUmC0wWmCwwWWCywG9JC9QHMx/N+av/3PBL//CTzOrbcRfLLRZlP1xcnp/f29vx2xr5/VCvj+v+sI6jtItzgJOrM+NUPp1my9sxX+SzfH6MThDsEijRsWhecYrg3jx1cr32ML35A77vm56aofNHOVh16+LiOtDmWcfzLE8dKT0XxCXpwI8AHZlFTx6y6IjBmdlkomQ4mCfyscPkHgFky+v7u7sCZJvUg4kMg+rBdhG0amXv1Pm75/7sn//vH7p1e+t3EpHzIaaLndk+DCBGuNDcAkBXgEfb1cnbAzzR8W0bCYzFIUSUzlOXijYCGKBZaQKgIR//gzlI42HdJSKU5L+2oqiUa7eVca04bGP/gdMFqLFcWoEIeXUfmW+Sp+WmPrdc3kuvLF2W+vSF9Uwtl+ful25DN07ArNtoHqnIj/AdzauzZ7ljKkAM8r766quJnju1vhFdAnLZDo5w2poZLy1Ly+5ZegGwUdQ02/KOKke2rtM8QkifWdEyARDMENoAB7QrH5My37z++vCPfumTw1MfeCprwjEMIl/rq57K4rpY1Ei9rhs5AcyKhnEtSEKb1mUo5HnkJvetbniFplghTS4CKo3c0wfQeBYAFAhbZfrwp/7Jl4Yf/Hs/wZpjgo2AiYzxAsAFTGgbVoIrRrs4nU85fAqOZVJv7DGbBHmToNVmynuIzl6rT/Xb4cDyf8PF8xvoxTMAUCW4ZxuZosc42GNcmdzt0iTgigqJFIscPLbe92YLPa48p5+Qu/PqWS+7xZbINNtnghWdnymUabF+aLPWN3KoEykyUCafbgfC5HvvYvyejRwTILuztTls3rkzvPb6K9iTpxQ2Alpd/93vfudwHsBS7gJATqd0HGS9MeyyyxRN743ezfiAUlt6KGP6eJRL+bRB53nvqzpjA9pKpXODX2gJffH0dZcNOXzPEiWrjMrse1fcUzoPE/PR65x8wVXHg+Xjc8mttupxKZBskmeMQJnRfzv8kcKdK12o36KmKT4j/VivbFZ5zXcWzLUc7aQOH9v31nzt4ms875bwG3m3nN14Rrr0FQnd4yNyh2v9CO/wwYIz46pJZvvAvMgGnXL8erzCDxsoOnUTuVxt8EwcHDJAls5++KPfPszzvj/c3Ubq3gO5Wyx7n9xNV5MFvnILTADZV26zqcZkgckCkwUmC0wWmCzwW9QCfDF3Gi8Phzu3bh9s7+2zyNDCFg7VAYAXfjDQAx/qrLWFj1vOkh/t9ffo+ng3ksGpL36t12c4jo4AAV6SE25qG8xa/F0yfS9cvgIAcHiLP4TyJ59THHCdOiNlTDoJcRTGSBckGJ2DalfHTmfMNaWKVrXwHpRDJ8Jrs7hJOTdxKGiMkjh0/qVe7MXyOCbASEYZHOCI6C9JL3CA84avfMCPpTX8wfXTp087/wk/ZZ7gEBpxizqRsoWV3XN3PzR8z//wvfdev3HzX4PHdzOV7uGKRAMEo1l2mNPGXBaQpVNr+zq8fVYWI1+kExTTeWyAwWmFRpJ59LQxIwucqmZS7mWArz1mcWZHRXQxaixRCfTD6QUigugQI8e0t0ln1wiH3Av6eMShTXHMqGwldxTnusr6osAS8cKSA3QFDTWu/cV4GfvPiJuAHQUspqzGlr1iGzVly/Y85uHjmMg98jInlWtE5Ly9szm8+LkXATOXs9MfGkcH5Qx7ALWADtz3pg2CO4kKtOVRp9giY4l2Rr3SQwJxEV/ZCigobWy/8qQLYDQCABXtgf3G9eEEGna2t4af+qmfwMZ7w0c/+m3DxqkzyKnN5Y+syCHAlqgldaZ/dMAFcBwf3ntddUZbQGekjoCXkST72k0dvKf5mFtetJ913SI/BZQ7dgSlHDdOvXXHSqPH5jfODZ97ZXv4337gbw9Hi+u8FgAPtTVPk8+F4PcBkY6gZDzrrpcESAU/U8bDeG3/Jpd7Lsfy0bAp8HoEAuyrEfg0SmzZheixJU8Ag6bGkuNSUN/1+toWMtVubHpB2wILaaarUKYR7Gv7DfkjoHYu+wUMyTgXwLByySevjB91gKl1HZf+q3FVCtV13jI2Y2nkURvHk+XaLG3DZ8HoP/Sx/c2t28Nr114bXnnlNfrsaLh+89qwRVSou8vu7G6nLeIeh7tZe+yJJ55IxKe6Co7J13XLavMTwCPWInSM2O8+cbanvfpQNq97zNs3kT36Iq3qofoCfWu+O5gqt1GWAoT9BxB5GHln3rx/jBBM4tp3U+rRrvdem/K80tbJud7TNmacsnyVVXrf45BWGi+0ve8+DyYT5jmRwPbsEqNDw9sb3jFemxzX6ZVjhmby22McB9lXhTbtz5ggtdCfe98RZuZn6yFl9DZXeR2TjA2fK4aN7dbvjmJU2vuOrD9QVC5co6d1Slbrmdfnzm/7ed9JGkxkYwDHvXbgIXtm0CcUYJPTvLMvfulLX1oDeN+i8w4BjhnW9S4tPnZ0JFcjn7jKnn5OFvgKLDABZF+BsSbSyQKTBSYLTBaYLDBZ4BvCAvkqro9y/U/2iDw83FxYXtxkQ0XWwl5Y2mLqn7gAURv+ldqv+Cjmh3tNE6oPdDMt7rMf6zriOlfm6wBlAfqwgEccijFiR7hE53QmyV8Q4IjG23FqB6LEKGdCJwES2FXb0pr6rEiphxNgKulzGbksQ0oKdIhOdJDC6Y1pa9gHh1GOcv7QiUaWlzmvHx4urOOQsM4YO37iWOuIyzPNEdHxse/43YuLq+tP79x+7ffiWH3L1q1bAFnDLjSCY1StSKCeste2Ohj1dkNL+ek0GmHitVMqdYDV3Xudp4p+sQ8FUZAbec0XbNolym8ZYE83SLvYNy7S77pGAVpwLs2fje5zR8K2s22oT85c5GweqWkkiBM30o3FaSv5lEtbU6zq2jblpYs52/vVTvWhdZTRxeDNbwDR/OhChJBtuZi6kXfu/Hfh3LmsraZtrSNwBHmmlHpP68dyd1vRBbdYoEZ5BQ5M2koanfjUJb901raOnbJB5Ukj4KItR92QXR5qSBblh8PNmzeHn/7E389aUufPn8ehZSfIka+6qpcyHB5QhymDuU5fls1jgzjcWbau5EKnKjV6r5xpcR7liioUlq51H53gaSodBXJ0sGmbcb4MaPf6nb3hL//V/334zJeuMqMQO9hRI5AqGLbPuJoDUBNANfoLzuHn1MnYarSBFTEf8mmfkimE/Gi7CTokIgkZDuDl1EnBkI2LGyHVBuohDnkIeKyz7zMpuGefZfxCUO8k+fL+oT3bRbMaQ8hu3wgOBRgZhYgt7EsOKHL2WTYpn8mySpWfMaJ+Y66n6Ay9Nbpejx/ls9+0Qvpkhl49b9++nfXzBK9doF9ax6/1reuz+uST7xruvXJ3xmYtxH8wbPN+dswEOMIWnvO8IId109YbrrEW+s8+b4nuQ2jXY7Qt+1Y72b73CwDOnn0mfI/7rAnEyNvr1sezNrDv/KMIIzdApO8Vx4jltm06Bub8WwKpbOfwKzrzmp/XWU8O/bSL+gkmO93T1HSx9Qw4Fl5jf2p3U0e0WTabun/7nD5kfIHHR2aGU2R0hMjLNk0l94leXb/zpWv5UoEfx2PH8YYc0s7Wa7rOt37TWRZ+jmGuZ/TIeqFZR/PoaAOg+57nn3/xCrQvwGef+Zd0CDV8/flzTEhXuhyP7y45setJznQ1WeCNFpgAsjfaY7qbLDBZYLLAZIHJApMF/iWxQH2c881MOMPB7h4A2QBARjSUjpS+jan8gWjsBzpQDEeBCWZKkGyuPcMoH+9+wB9PgZNmdApkrHMlPJIPfuokCmeMMJJHDhyS8qmOv+lD346BDls++Wm385TH/OgVoVTCXGggNnpA5ikfHSWzykcowpPIpYpSULhM7bK5uaV5/iS/sjS/tLp3dLi8c7CHd6+e3eY8nrA2ml9/4sl3vI+/5H8H04Ie32IRfcEL/qqfKTHS6PDpyLcjvLqyTr2jREA5/aoX594mSmQFMGIbcOyQ6CCnDAqEGVkmSKD94zwCRggIteOsTXQo3Q1T5/uAAEHbMkLs1KlTTL2sqVGWLQGiubtjmUTAwv5pZ3B05rBbwIXYVYtqN2wWhxn9Rwc4eWNZjRftAVlI4eE/jF7Tb2mDtpLS77SKnRM9CO/Iy1k9gAzS/9rI6Il2NkUdX2dR8xe/+MLwTe95D2vJs7Yau/85PS2bAlS3pq5RVmhZ7SkTB9XRA+c9jjBrW5URiMQq8GVeZxkaI99aNxk0MOs4pkQzhI/6OcaAEzLmXNReWXbpv5/9mZ8ebm/eIXrsI/SvO4hKhZMNsKTjbz8asVPtjP3q4use6Gyy34vO/qKftD/taxe7xoX0FVjdrSNwJOjRwJ91wwdaQS+jzhIJ5NTKtY3htTuHw//6f/yt4bkvMmUVswh2x1DwjVzwNMLmiHFpO7WY+AgUHI+BEUwSWbNDE9XmGFEWwEvlVdgYTWkoS/AlYw8eAiDr6+tEs7l7K2stsTYXqHXa015Otcu7gz5aBEjMOMmYoq00XX1gz9BR8LQ5x1r1YcCaEfiwbU1xEOCt5FYiAXr/uV6fU8QVVZnhYjGq1/sr9ck3N+88r9VtPGsz780yeV/9cpjplQJkTrM0//r16wGnpF9mHTb1uueee4YPPPX0cO7s2QLBfG9gI99Jm5tbwzZH+oX6dCdJWQGwsJ3v2az3h1FOop+0g+JRlmfe58RIM2Qc1+mTS4FkRUfv5h2ifv2u7eg4n2tTdOQmI5oGslsp+XnvjjZQbqfC+mx5nX7ALj5/WtAIVpP6GJmYsYqegn/+wcX3nVPoA7Yji1FusXnGvBz8B690O3oij2Nffj6NnmOrtFIyj5fhY5lArGfljq4OHpJrDtquTdUgO3m+8gch6sBRpo669EG3pW2iu2Whqzbk5H1sN9KYZ/KxkR2TKEseGpYWas5pxnuqoiBJ/thrdW/u6D7A9/sOd3Zf5UV5xxb4XyODhyDvOvlbKT+8kN+vla1Kpp+TBX6tBSaA7NfaZMqZLDBZYLLAZIHJApMFvvEtwOdxO4QHBzgDd/hI3kStAz+Wf73UH/OeTXV+88c/jgT1dQL9q3aiCKBdMLIDJ9apRaIRsjBKBjdOTjms1213G7OimNf5Og8ByeK5Up2UurDy7FSq8Kui43Lrmy9YUgkgjgvXVmreltd1nzEK+uBEosXC8u7B7qr7QbLmiwLTFE6K3uUw79piw7f93j9w+YH7H/qOl1+/9h2bWzuXcaWzuPj+3u4K/gwYgGDZ2DqOj46wZsk0N67ZOTPASTuj+7tw2NuO03oMcOgqIacgiXQ68cosL5N05u8TdRNHFIc+U+poN/fQCI7FRvDpc9YSwiK4grQAxNCCanCSdCZ51PWoyFhmsXLYdtvQqDS5+V9gyXqzNMVHhzkEKY9NxjbaCbddaS3bA0TEkji0h8NLL72UKLvLd92VjQmksU7OXHeKPfWASbbf8tU1vXcsM3W70sy5y6te8SjZi17ns+wXfzQ1Q0tb24AgP/uz/2B4/Ml3DJfvJhrIfsb+mfZ4LEvx1LYHOxVBZj/ab57l1XZpsZRJ+uhGZvoWukRRxc7VT7MyS6tZlD0AAtM8l4gc+4e/+tnh//qhjw+fe/XWsD23jG2J0hK4Dp20GFWQiz4M2AXYatRYnjUi/ezg8EQeU0WRVr5riUVWxhSKBLSSL5fhn0g0762XurX21KHTnMl0x0vBD4GhvFvQwfb0/R2jAr8+Q++3i4cAACAASURBVMpY7ci7x6hNyrmSMnakmPn7vqso8toyz+AhbwA5rFnl2g5bjLqKZAhIlU1rbKcPqqnQ2mfWMSm/4NPuTSJKAT5Nlt++eT1jZJmNNXwPCJDZi08++eRw6dKFY7DIceBOtXcYT0aUzo4L23D8CXYJegnoyFvZ0o5y86ryrmiNHhNkQgYANZ/RY/q8VwusNJJM8aP3qEddQz/eyz9YTfreKK/SVzpKMi6drm/3E5cGMG1e2dq6WDs/K6LQfoA3Mq3OrQyXsJd6GtW8L2ALbeRnaCmz7ynrOVazaD91CzYKy9Dad51Kpr6r85vL+17xc011z53ftd/8/MpbmvqjSsnpvfldNnvvWDG/z/K13CNjCtvZJ4556WbLuRfxSibk0qyurK0+QCTgg/wCeYaX5B0qVceN8ocBPxzBs8n2pjRZ4Mu1wASQfbmWmugmC0wWmCwwWWCywGSBbxQL+DU8fiHHHT0AcNheW1zYyqf96OBCk69mP8z78EPaa89+tMfj4acf8eb5UW++1+bpEIW+/J+UJ6DE6AWcy4W5mlo2fvunnvTyqbasWA53RQTAE49Zp07H3IiFLu+/jlu/JC9nI/dQedYRKQcW/rGAPE6cElW3ulFMOtyxDj8FBfDn8IXnmEk0v0T5/MbGhhwwyLIeDdeLwxPv/+Dwu37PH7zv+o3b74fXe3DcFvZYLAjwZ54pXotEnmRhfmXQTupptNjhEs4dqiyy8+XqKkub0Z6RJZZvglsuHywnkkJA0Yivo0OwOMrUqYJ85gOkIE9AC6dWxn44l7blNFdBhKX9AsUEZ7ThSdLe9mvJpP2srzESLaOVtB95tqndBUlcJD90I6MCKGpUSKeTT0XqVH+etFdXBaDWcFRX20238MP7faKFlEv7e8/oijxG9ggEbG1uDy8+/3xkOnPmTGjstTj6xbb4GAkCOJEQERshRT5s49k1zWBMSbWj/bXbLDhnHWVQXwGovjbfiBrYJEJGJQIEJnqsdq/81C/8zPCFFz4//OF//T8eTp05Sz8v0yfIQRua2aQcyr7vGlNc2s4efWbfjeLlWvjUdecWiLhpICxV5SGjkZ+XymhqwCDPJPc+NWid9cUW2LHy2S+8NnzfX/uBYXNYG3YXVhlbTuOkrt0Xrjw3DjT7/AjgzDlojPesb0TjAmAaoHdJzJjgQT8GqbQZdQmihLfK+XDBD1y51lSD1n+0p367lFVz2JudI3cBepdU0jqkGnPWIJJS8BBZ7bvC8xx3TVfvInUp+5ZNXPjf/q015OjrsUbsoj5WRxbHZ6bqCrbFXrbtWLGcFhGpbCxIaW2izthRV/nSHroGmNaGCGe+z70RpQ18Snf16tXwsX+89/k8S9TYk48/FsB8+85mnv/bjPdNALID7OGU1OgAT+mt63OhfQXhVlYA2aJIvZ+NEpU3lkDOGd3QMYCaoJTvbORUrwBeajTqkmcb/dTXa3U1Kk+edWAL2tA+Rj5ZnneENNJCFzt7z2GPjaJQVjJSicQfFLBtoDyeoTX+HGE6N3c65+4zp1/uu/Ya/ejzYT0jQH1f0etpz+c38mOTnCO2z6/9xfgOvZmVolbfcFZeZfR3le88dYhN4dd/ZEleCUCNk3EmHf9TRxpTZBh5zF5bZl/GRp7RO88L+ebZL93XaU/GFnEI0HoBP1bm379nZ3frHl6cq+nH0g+j9JtsbIP68ml9Tywg2ylNFviNLTABZL+xfabSyQKTBSYLTBaYLDBZ4BvTAjPfxJkkwgL981t8hCeCrD/U/Q73Q95kXic/1k2W6Wg02OM5H97Q9ge/NCd0Oso4J1R3mp1rTOmGONXOiDI+5POx33XTCE6HNJ1sz8ghP+5LphO5vCp5T/Ks1zI0jwJ9bJsySLu91tsdIs1bJHqCE3NZjub293c52L8PT1jA66FHHl6cX91YPtzb28Kb33n8fU8P//5/+Mfvu3rz1lNEPDyGA7WwiyNs9MMedmnbGPnRNlMugTCnPdq2+Tq7ygQAl7JVokqUJc7zUGsNeW3dtnv0GO91jk2WSSPf1IWnZcvLKwHlzJ89bFvH1zwhLu9FLDwLjJl0xkzemS9QI/2sfQ3SgnPVU+5ErYw0qV3OsDrJNu3Ic5R1JMnJPOlED71WJ1PVYVwRYfTpT396OHfh4nDm3Hni+5YSgRMifpQu41nZR/nVQn4muPKzxqugo/lO9VNXwQZdy94N0TJ5YqnYwPret60dUUazaLrQcbHNGnIf//G/x2Lrdw1vf/vjNaZGR7qn5y4u0T5iOFbkhVUjxx5TGb0XEHFclM3KJpFTefhn8l657CvHT8taZdVPLhJv6sgXI32WVzeGH/rxHxqu76A7u9/tM+Yz/RK9j1aQAxnEhEBkUremuKEpAjvdlQsOWjaLy9gcGRAgRxb5lwynPwCl+dh1jsg1kTv1s07+McX08HB+uHWbacnUWXTjCBgnsoixSc28KyBPHe1hm2FpR9kXjkn+xR4OYYBRAQeTeekrOKXf7OdxbHW5Z+34z0rpV8oXeHfJy742iDQ6RQRaV0CSIEqeH5SRNu8C+tKz7wGfR8+uT5d3AM/12toaU0w3hrc98shw6eLF9LkRiNvbu+x2uX0slm0YbSZ/x0bO6Jnp2eRFTs52ecsTvXh3+j4wCWYZ3WsfWpZnocyY8qbRvtnQgTaNDMzzJ4g18rEfgg+OdpNvntuZ+5bB/JbN/jD53gk4Lz1jw8g0N345zo+RAfJ8t6Gj43sJPGhvQZDQXS7ZzMK1I5EpwBI8ine9h5Qn42FEiivSrGkiwvGPyDl2f2/+clzIhbrbrz6v3acC4vI/0eekRueZ0zY4KT256jLP/b6lQniWLavtbgc55nhPZQ0y30iAk6uUXXnve9975ZF3PLHy2X/6Kzy3KHI8j73aank8j2qeCDFdTRb4MiwwAWRfhpEmkskCkwUmC0wWmCwwWeAb2gJ4b4db+A7bfDTj/xSwwjXAEB/hfEjHIUJFr3UKOhndo4NitIHndjb5rh8dhnJQ9LCNeHAmYsAdHQx47XEYfaPjo9Ouk5a/2uvs2i78u23cJvL8rzw4oXh+hzjtliuXB0zrXiruBdE8y7McD4SEpgCmctQgyH07IaFHvnZYXEOq3Gv8L6LA0J8osrn5jTMXFv/4n/zTyz//c5/cevDhtw8f+/Zvv/DyK699BKfk2wHW7tneqcWzAcfmid6KHXshdadJKYO29Gw0ie3q3Ors2rZO9IpTrXDw90YHWJp9dqYUvHEqpuvzHO2i2xgdEucTewqoyFc629BRMlJnmeg0puFAD+gAGGHERZxRd4gDnLQfbCNAGO1mvSm9UcyGUOkdfS4tihlDG3slT4fRkQEd/Vd8ip99pjzpWyjULf2qcy5/nPa0SZnnrGGEPKbQ0d8VBVdjb3HFOKO54QvXrmWK5dsff3xYO7URWtfFso7t6fAjJuyxGfdOp3OcKo+6zSYjhWi8xAEg1X3MFD7oXBvMlGE5gohHeMhaJCmONzoWSoBdG7BYHH7hl395+Kc4q3/03/2jwzk2EtgnIsoIMse7rXTEizYwpY/pj/StfYFcHq5B566GJvtZOv5r7jHZXzxBAgiUx94qa8LGjoM1ADDbe/3a9WF941QAFuOvXrrOckVrZ1ion+l0jIF5jljAd0E6XD70lfbhH4MyfZxprgAmFGjUStjLPoyM5HhGGC8CbmQ6HH2U8SE/wQv0myMqTZsuzC0Nt27dHG7c3BkurZe+0jotMsAltPu0r63DexwnNk4rSdKbbDJAHNdlL23GQR9at95bgFyhhhbeVV7P/8gmz2PeB2mLMmzMG40dJ3UVkd33jh1x3BcjR8Twvee6aT7jTMumXRbZ394MoCOXG9deDxi0CNjl2nQCZWcYy48++ijsFgBYdznczZS1wNDZfrFvXadtjSgxk7qY57vKs6nfX+pTzwO2hs570R3zBHYEvKyT5wFZTYnyow+1h4PePvP3grfFFx7jHymkt7/zrkW2slO9Qw74A0HKE1lWfZKplsmFlvaltx9Ch/2Kyo6TV62V2Lq4Vp9/WAkNepjvTq+CgIRBB7hyPPm8oyiCjWME5ulry6hjkXZQ5rQ79nvxw5YwTLmF4RPFaVdwrMaVz1N2EFbnkU/xVq7Sh6aOU+zOnTSzKe2MeU3ju61SMe46lnv4nrb9gIHAZEsLhmbaSXPnH3n4bRf+1v/zd1a+/y//peF//t6/iLAy9239axOWR/o3FrUOv5Z6ypksUBaYALJpJEwWmCwwWWCywGSByQL/slng+IvYT2e+t12DbAu3ahOXad+Pb6d2xWlyjgypP8z9eI5jxVmnTN/BZP7Jh7VOUTn1mR4nTdrBcYDdPo6+i0eb5GXESDt4+FHUJOHQB2TxMo2UQ9ttk5v8gCmjELbffkXLUnVDPfIpWQ9xsAU78HTLYbGq9WFgG/5DpvrrvGEMJO+JmFmB5ylss7a1tbP60W//nctPf/OHiXjZGl569erbd/cOfjtO029j7a/zO3tOEhNcWVik7hERaPAogFG5GhTT0TFaTHBMGfpQjgbLxJAElewT6x0wJdNz9EQ2wSMBlbJnOaXSsv1CaIw00cZGoxmhYpmpdK5+CC/k0tG3D1S6+WUnT/sbUwhsdv4xD/KObc01N6VHn+XnNQ5xp24vUVqxfZVIF6eNs9ModYpNyR/52XfLq4vDK6++PGyz0PmlS5cBdVzXayXOo/J1e7bjKM597Guv6DIWX3kXjZ5vgQ/m/XopMiPPkevnwUsW2tX2vDd5LU4mWHEI0PUjP/p3ho2zZ4Z3vvPdlpJfa49ZT0nCB5BC4MRNGOYA0KqsZA5P+Ak+S+t4WWIzAqMSo6fajGZNn8O3ZQlvhJR2h0i2O3fusNvnWcbaEuAr0/A4ltcXhgt3XRmGqzvUYwwi397BdgC8DALHiutljQCe8iRyDJ6JztKMc8BsABQ+KVl7DL7aG0r6XMCX60wNxnZ2nmWATeqpzII+0hvZsweosoUt7tzZGu5m2uzhaNvgcLG540/+Ambao3Z+TH145Tz2v7KazOuj7F1293k0KUfbijuuqz8zvRJ5lauS9SjLbdEoh33a9W3H5Fm+guKO4V0AJp9h8wVWPAuUv/LKKwEqBU19B/j+dZdTpwzvssmG/V08fae6kUeBr9KtEDGZxHOFypFB+X3vWsepkwJ5SIMs9EV0Y7CkC0pO60ub9wv9pB6dZ59TBEt+2Ie+Hew/8nMyx4bzXFteqW3R7xnrlg49Nul7GAvYmcLCH6Y02LqUbJUtj6JHKuQUbKw2i7e0J/3YMli3dfL6zanp3nBOM9iw+Y92az62Z996mLz38I89scfYiHnNd8wKXdfxLH3z8b7b8Lrb8dk3WaZNs2PxSMh4xJRA+UV0Do7nAblXv+l9T6WO1friyznb5pQmC/xGFpgAst/IOlPZZIHJApMFJgtMFpgs8I1qgXwFj9/CrOu7v4kPs7m4uHBwuL3VOvndTRDBCDbwca4T1cnv86xBM2aUYyBYMEaJ4VSMQBMU5Tjk45tG+xtcx8A8eelYH+Bosdcj0SFZ8YXpVUXLH8njGOjrZR2jsU4AOOqWUwgf6gf4GEEVRYsfwZ/9Petseo6stFGONvWQVT+C1gIClS5IrcNlvjtQgtYQfeMCYWcBEC8sLC6eYs/Ppb3926du3t68jBP8ASKNntrZ27//9u1N19FheaT9OZYgY2O+hcAL6qsMuyw4bVoiAmTj9EaAMCNCdDR1/hbxwHWAvRccWz50Z0bXFVoJMCYYtreHnbdZYB3wa2uHXQWx8SFAhvUxYnQsu6Ibra+z1tTG+qkc5r/xMMjHiDOHhX1YQIOOcdsiU+XogOwUakRWrFZTUY30yz9klYM9YrmOsd2TSBTzubG/8SNJjg8iRKyAnqbjtuBnxJAAqLsZVuQXDikgwyKgQNvimWeeGeYADFyvyR3uGlCUV/SjBZ1cZcjYS779TRQXmUYw2rwAzeie13iUwkqc47xyHdmRc55IPMFO+QkSGIHnmLM8wCvnRXYJ1dY/9ZN/f/jUp35h+AN/8DuHe+59ADvQpwGGKmLQSMgkukiQM4BvRkrJPw/QpPACHUlG3JH6mfE6USzoaP+1o+119KXeHmPlNlP0NtlB89rrVxO99ND998VW2nGLR/ouNjhY/PQXByb/xhbDEe3yPCqvO/ilw8aonDnkdM0xwQ0Bb3d+FTBi9A2HADrK6yj0nATd4QFRaY4Z7HLgmKKCgS0daSOdIJpNKBP4HDuTfml4/P5z8K4xKLC2T7uOlVpryjHICwFd1Tf9Qz+YnJ5n6j5PXyWjxlX6fIxusl4ioCKPJb5/SnxGD0zIAqjldcFp7Af0q3oSluyq2/rwzLNBhgCKwPbBsLW9k+deQMc/PvgOEOD+0he+MLiT5ZV76A/eBb4DBLFPnzmVjSdeP3w9upln5NX8/Ar3nnl39ZlrowID5owycIrYgmNtg/6jhPeOf1OXgfx7w2HfcaZ/1M8OsT2vA/5QB41TX3ucAIdUJUPrGBfpdMx+lsnK86GNI1RoyuYlCxmUea29bEtSeY1/myAfqSgcuyy8pavNFrRHHQ26jt0fPrAhOU59Rk9+l9V96eZ1H+ELfcmBIHlBcSpG6bsGLa1jkq8yn9wXdY+HY8VHHvJuWs/ezyb/aGA+b+TY/Zi3ckKobX1nyRdgneC/uUMeAXN4HS6dYR3DUzdvsvurvzze3Lg56UXfwBh8JrUUpdVMwXQ5WWDGAvx2mNJkgckCkwUmC0wWmCwwWeBfagscADzcxpe+zYf3nh/rcVIrdKejqOIYjPn5QBcsk9ajnSHP0ui8ZSoV399x3P2w5+BH+GjNWXBMZ9EEQEc+n+mL0pMxOgoCBA1uHRFxlg94HGZaST1lMNlGHI7xuvM8217T9bXnBhNaF50xMQGUGgEAnJAxlABap1ien5tfuA+KK9R5+XBu/gJtvg+9P8p6Yg/vMrVSWI31o+Z1+JYWAbVcVB/ZXG/INk22Z9tGdxkx4jlTLF2bqctRq9cZMq+n3QkEyQsOOctbG3Z02O4uEUC0Y76p+odd4XS0adM+8tz2aBpcztD3D8sD/hjZlMz62eWepbGZaqvGg93RY6LbKLqSR9rOTz2y31A+2kgelhslZP+rU+tl/nPPPRc9rly5EsBHu6jbG3gj40l7o+OLNvLR2d+HT2QQ6+DadFJfQHUcb+T3GAzR+EM+tumwDQgw5p89e3r4kb/7w0QO7Qzf/tu/AyCTNZP2aGvULW1Cm+lsnNXVtc7kZ5oF+4xGk14aD3GhQwap8tg2halnn3aSzqilazeuD1evXx9ee+21YfP2reHUWkUqSuszvE8Vd0qUz9auIATt+IQBjhmlc3QIfzoUMBjWtCNIpZ0Aw4woFEAACiaLcmnsfEA0BI0omT7pGJnnfbHPc06klKn7W3WdIuwjJjC7Z10A7hdfehnA6Mlh90aDfwLHJ66Z9R2bbXPtY+8ppXliA8UTu9KI/SyQ6/NNLOhx+11PkMkoLjkIzKjGAjaIvX3XmKFZ0Mvrlt9zaKwJb/uk+9Zrn8vu031s1M/wzZs3hldffXWMHhP8doOO1bwDTm+cDUCmeX0nmBwPq+P1POMh7Y6Aj+Xe26e25XWivJC1xuyJvtKajum8tu9Moy491uRTh5ZVz3qfU0HSJGl9D9FQngHpZstad4mzlpxgHCk2GvsMYdJOWhnbDBE/qv2SrwCzGleW5/cCY3SXxfrl10cDU2lj5CG997HNmDe+1qvtN5T5HI02sSKpedvX6qRd1bXz5WvZbBtemyxrOu873+uuY15f5488FpLMLxsUDzKqgJ+dX2T1DsCSZ0+trZ1zqi4E9kaaPq40XUwW+CotcPIW/ioZTdUnC0wWmCwwWWCywGSByQK/+RZoZ6IdoEigJxlfBDdL12jvxs1rNx6eG64tLy7u5K/xfITnr/ZQ9Ue4zld/rBMS5Zc7EV5GG+mYlXNg5Jcf+ZkqppM5Ogzz0FrXaIrwSURXywar0TCusyM/sTmBsjgMTt8CDNCBZweBOHNGruD9plY7H3VWXpzC7KCHw9EOjM6ch/VI2W1NR5h/6mmyfp9ripIOcunMBEl9VXSIfmdR5SGi1d62tLB4mwCnDWJYPrq/v/P03t7+OfVURw4wBaLFALK2WcdfR1lAIt4Kep4+fXo4z8LyRu+cZQqejnDvPtkWifzIaL5O2bwL7LMumc6ZZUssqK7j7EL/ph2mbDmt74g8aZxiqSw6XNpPp2kNHt2P2tfy+SXBGaaq2a+kLlfnRPsYFaJ9ylSJ6gnQgz0q86QvrG8fmsqhDZfRvgXaGZkUB53qZfdy7pQl9kldHe067LdebF2Z1e2ll14avvSlL2Txe0FE12RbJkLJseh6XSVvjTGjZ+xn82w3oN/Y30brmU8YJYLbMG0FIVUH20d+gJVoVKMgkWOYVEPxQwsAtMLHPvFYBQx79tlnh0984ieHb/3W3za8+93vHm7eqD5yDJjUtWS0b7A7NtveE/QcAEoKRNIW/UxZx3tlz1g4cC2u4mVZtV2ggTI7rB0Xn/3M54dN+AoAdYSS0/pOM+ZWT51jB9UBG94dux0dME2XNcBMi4yh9LHgBd1r20aB5aaBMPpBY8RElKdRd7nUto4lUSqXR4JmgTXGHGMLTrWEVt1d6N6RY+Rd1grjmXbjjiP687VrN1MWO2GOLfrH3QSta1OxBdbKv+oGccOk7mvpfKfUu8xeIgORrGviDRY5HOPuCqr8FZlVYFONHvt27CvVR9n0G/XdGdJkxFrJVX3j+NzbK0BX4NCW07HQOs31NkDl5z//+SzOfxZw3GfT3S9d606QO7bBfgF8GReZCks04RJHtY2dMmZ9X2bQRg53FY1EpWaeGZSibARX1I96sR39avRjrkedfF9535s5OGbmGA8Zn3DJ+zj6+G6lXWgjD/USvQvPk1S28D7jNbYre6UPlIUL69umeXRDbOW0VPM9+h0lWGub0npQVP1K//JUs9YbUXv83kgdB+RM8n3eHZC2vJM/wH/eQ9zDNfJYTb1NAQ5hFb1p5Qj+9q3iyq95WS4/k9ezqWk6T7qSv+jT/ljXa5MAtXRGiXUf+R4wgs62lTX5sJCXzXv2gMc6v2su8keX02TcIrcfixaB82w/zWRPl5MFvgwLTADZl2GkiWSywGSByQKTBSYLTBb4hrJAew+4rbk82NveeQ0n8ot8aL8K6PMkYE8+9HUG+sNfDf347w96HVcKk+e1Zcs41YIjOh5+hON2xqGQh/Wky4d8ADC/283HDdAZiOPhBz5OCI4wS6vYZNrXKbWe4ALNlDMvQIb4b3ZIbMfDJJhguXqmXfLLQUlx8lMOnckynbbICa11zO4f3kO/zulhgKj3EvEyf3pjY/3mzc13bG1t38M0v6WDg93DPVZi12/T0dsxogw2rjdkfZ3eczjFLth++fLlTA9cZfF8fTrLlaHtLtjX+rWclnWei39bR7u4i9v+XjnVSt06xBbQuCOn4FicbhxyedSBDQUm7M8xNX95eyBUSsp2cj9JsZmdQipHtMjNf3MkR/NTJq8929bx2kJj/zT37kd16SmIKWN8CTC8/vrrwze//wPDOovPtz7yrbaVuZzR6EBvC9j6z4g0wc62uRFFVU891K+cc8GV4nVim/DSJjNJGpNn5RDI+Jt/829mOuN3fud3ZqF16wkQN6333c9Vt8Z11lFjjNinOsXSpU2InIac0TzWdaqhPFIfMNdUPKnD2LG/77333uHlq68ByJ4abrE4vwDNOaLbBGyXsbc2zg6A6a/SQ0gnIDf85gFkD3c28xBIBwqRdmI83iDK43OW6DEhKk3jvX55piTyLCJLxq27wvqcD4BdjEH1Sh9j9gDgTj323UG9zz3/QkE7RFQeADaZ2haz1p+15+z1LL3Xlp2MN3Mqz/w+BP8EqTArep3kzz4P3YbngF/qirwtm/m80nIfUJw+M/VOtr4fHbcvvvh88p367HpjAmPyOHPmXJ5dC1cAE09trAcU97ntBfWrba1Q7znlExQ2Iqrlk5fl6VGvabdlrDLH08nzZ54RWdbvo9fUmuVplJ9gVWhowXP4CXj1ePWFN5Z51paOC0alt6I5ADzkUrcTrWo0JHZMwXMskHc/J0xyF9I8btNdbAX1fFak83gDz5bNNse2msazSZktyzjsRkd685uvtN47pbnlMa/5dHnTS9uHZZ1m6Wfzuq3qk7FdCBSJrjvuK8tjK8vQwXej8pi8pnztaGH5MuD4ZbJE5S1sQ3ue0ZK7KU0W+AotMAFkX6HBJvLJApMFJgtMFpgsMFngt4IF8PB+vfTGT2PxAQiPDp5//nNbH/zWj7xIBMILC4tzN5ePls5s7+zin+ug18e6jl1NQ2INJnjLynWcpHHKjw4c4NqxU+AOZP0Br6MWQEIHQ4AH4EyH7sA1s+RPZIqLcUuvA6ATYrQIxOGvmLZdDkD99VwBcIeoD/dEF5SzY6QRxKU97cnPAAJ564SYsg4S+rTj0flxPqDRAUQl6qS+8SOph66wOVJtVjU/ejfrY62ePr2+f+7cmdM3rt862D/Y1RmZx2Gb297etT1ZzO1tE51FJMbS2mIAsUsXLgznzpyNY2zkmDapqKaSWz2V1+S5naB25nS8q28KcBNcWF5iCt8StEZfGGqgdZy6xtUy/GxndXU99Yw+8MDkJ4l2pLW9fcDJtKXhxjyUOfayqi/oXyMqbIeKZcOihzSpplQpowAJ4IquL2VtZzsv9/a3/U9fpZ0Zwbr/qu9ZzJ4KIJCs3/RFQua2htMACG5yIMDgFDkBjuy8CJ28IxcXmU4lcjGCjuqZtX4yXMrGThlUZetQjLhlv1GdyK9djTBL/0T+KrVOIoEYOJ957tnhR3/kB4ennnpqcLFsgVIHgpFIXJWN1RmOcW7pJ23oFLuyIzI4AEkCxspcGi+1JAAAIABJREFUNz4HTBek/xdZs8o5vNLDGQARQA1R0m/2pM8LPC5dZMH38+eG6zevDS8TUXb50vmsj+Zabv8/e+8e69l13fede2fuY+48SQ6Hb1GyRIqyZMmKg1Rx4jSJ5KKGjQao07RKUaBIGrRAi7ZIC6QPpGiTPwK0/xVF0tYN6iBJXdiJncSO7dhxLceKbZmyFCp6UnyIb3L4GnJe9337+XzXWb/fmQllS8ofldizyfPbZ++99nrtfc6cte7ae6vbRNuhl3UimFwOLFdO8DiXXe6bMXE+8tRHKePcAoZ9+NiqzHEl2UbdsIhqw2Gnvl1+pwzejskTRXWMZ38rZR+de/LuPnrMiuH5558frnC45nFO1jw8dA8v55ncOSZLp4koM5aOZ/ijgnFzVLpenS/mKO8H+5vizFd/XB7yoEO3nr1i1mekxqP0fxyHYCfxy01wQTfzlDF2PH0+XUrpEld5sC3POPk2TsCvPfHkcA1HpfPU5/K2226LA/gE90aSneCE0Q3G1zntO7X2AZO289JnZnzvhj/xj5FjlH02nWsmuTO6LRvr+2ihF3lRLnOTuXr3Ui2tQ2n43ssVOq0LexV+n+/Szzi49I/mfbGSGhdAgWve5cx+Oa1WuAJO3zjO1umPDPJmnzwjI87wOcJnXzr+SJAEL27Zl0Tf0AaN0YHBT0PzYyCkPDmXTAu+oOW98A0bgLHsvzO0pMr20mXNjcZhLo/mXdc4SlddujFv+JZPWP6MAY5yqlv25NvojedJOOcr7weq+gURJ9k6f6C6/eDw8DwUXuTSSSbTkXq8J5umUQZm9JxmDfxeGqjZ8ntBze2zBmYNzBqYNTBrYNbArIHvPA3EOtBY/bVP/Mpw9fLll/b2dp7EQHyej/U9jGvsKBr5uOZjnA/s0RjXsODjXEOyLx0D1tVHe7Wrji77Ud/36cO6RPO19XLcmK9vHGdZF8Y5l862picejYfOvY/dnZr6sa4jNLy/+WpDK30xumJkiGc0EsUy5dF7+TPvC1j8N7gN6Icsm9Tfz2blH8J8e/ett5xdO3vu9FWW63ngwcoefjIM+sOr17fNs8+QG8nfceGu4XaM4Ts5NfDW287lRLrDMfpBHprPRIRhaDe/HSHRxnfzpN7l07yu1cU+Rhre9rfevBxky0gr+5kcl2mkkrhN9jFlVR11lrsu9WN7gBY/GlhlZDUec/v1+Dfv3d5topjWdT9z5U4b0UWtiy994fMx+4yQ0hGknML0mEqvk46I9O+KMZf2tL7la9GmOG7qutBH+o9z3/46637ll39hePH5Z4Y//af/dJwc9hWXTif5a2eJsnRbHMzMe8dF2L4sT6+ud5mxePqStvuHFf7ROGcIO7ru+WefSxTjm0SRufSydSo+N4A/s8XcYEpYlk/TQpfjXEHoOBbSODpbfISig4ahPxUBiVfKPsjJyOSQBQ1+nXdQCX7p6UCTlg5LZbX3G6+9Mbz08mUse5gy2g8Y9RU4cE7HbaET6Hpv23Isl++DyIOnLH3HKKjWt3XhBdouaV6Dj8Ylr+GbtindErL0ZL34s0G/fMK5PFRdHcrgBv1PPvnk8NTTT6bevQd1jgnn/DWi1DqXbvq86vaQh8YjPe/78lnzvuu73DqyfvkULPumAz83y2LZeWhu1G7GgvumMe037Vvwy3flzXANqyx9jT68hUO6cTQtZa9+1cc/fHhIx81zwGXVOjdbT92/eTBv+k2j64RtXU37CTctNy5e/0WfCXpze/cxF2enKdxbtVln6nx6333N+145he0yOYGxusZHHEerBIYeXuAE1AsA1gZ2NtZUKGJVnn9nDXxLGmg/9LfUee40a2DWwKyBWQOzBmYNzBr4/0YDyw/0oj81k6xJuz/YISvDz/zdnxpefuX1K3/tr/+fj60crDzOnk13Yx9lMyI+xjkhy4/+CvPw4z/GC537VDf/6u/VRuTSQLjx4x/XAN/sGpT9V/YyNI65BxZ4j2OYxnmA9XRwgME6Gg9l+JXDyD+WZ2PzMAFcjJE26F2CqURlQIhTQ8I608IIgb4GqUmYZbtOMY3SMpxsF86IEJyFHFiwvxJHDPrDgDxB3T0cb3ny2Obq6+fPn9u/9PqbB6+/cZkIJwxlnGObLJ/ydLo1HDvuK5V9x249w0bpW/BdSy9DfxIt4R5M0yT/0UnkLDkwl5CrjGfb5F++tog42VllHysGzwiWg4NxvyflIbJnY6NOemzDVzrqZG+MAnIPsjK+KiLEiAnL6sSR9F5+c7ph65Xy/grwAJTRVgZt4V46MmTfkSkYW4EHv44EzNuRjlSKjnfyGfmQJ/sjOeYYytd2LrNB/1eHNU79u+OuO1UEFzoxwiP8SsfLYo2luDLrQ6HGPUxTli8jmpzh+DPRZTkldAvXvB47Qds5yUyMHDoWo3ty8fs8vPraa8Pf+ZmfGt7/wfcPP/RDPzRcvPhaZOPQBozrOE6LXVHyXLkcczEXIe58VnYjX5qOS/9qHJy30MrzQau+JmCNeNSJ5NgcjvNHB0+FTTE+nHIqjbvvvIvosY3hpZdeGu4i0m7z1Ik4HTbps8/ptfvsl+cSR8fbnx6r5EQ2Dfu8EpwrOLKM9vNSfiOYouxs7D/2Q1eLJEKeOYjRH12vcOoqMniKrDybCA5L9JTt6n2fCMxnn3tpuPPce0q3yLPCSaXOB11o6kPalnnCU9bRZ1n+Mm+AdB7AUWSJXAzyGg76VXDpdAseIJwDx+FnDf3CKCV1rhpUhnPUvFLNKegy3p2Uw2XAviukvUuU4x7RTTWGNZefe+7J4eGHH2ZOXIwj7N533BeH6jGWsTp/zp0+w5Q4Yg87DuzAUeX7VBJZsg4fifYj1+mu7AxVErfoUR6jGeSv9yzSoTMafRBIgruvYvZMC756j3SkXO+56Jz0ne+45xTRnGrKAFGn7FAe9Sne0q34TTVPfZ7Gcc1DONbDS3CCw2WW1IY3isvk3KItrfDou/iIfws87EGUOcgCaPW1Bqz0/HdFJ3jGHpz2NlrO/+TDfzPUV/CCO8+0Yw+RQGUeskzTIeYSp/iLV3Go35JHgIz6yCfANAZR9R8leSs9iK/5aIHF23X2EUadmiowTBlTRCbVVe8Ca5onpOfvXHJl/2GDE1RvZ95fADHhydU3jY14UdU3LVuX53zWwNfXgO+ROc0amDUwa2DWwKyBWQOzBt5WGvBDnMRX+CrLAjEM2BPok7/+icvPPPX0I9hPn8GYfskPbo0hDCVsL02qcja10eB+NdMPfo05P/SDOB/5fsxjhIwf/TFUJEqdV3/cC69xOvIUHCzzTESZ+LzkpfgZLQU7kd4Kl3XT1MZHw3ebxpSX8NKe0m+8zXv3tUwfCcSiQAZ8iQdnV4b9W245d/rkubMns7+1zi/2GFvRIcbqS04JPJ9IEaLMcFT0Bvpl4KgHoyKaH5cP9r3GtqdVmt982U9nSpbCoSMjP3SC6IhTV8ptnbl8b22eqPrR8FUE2zot9bY0lrov3cFRkK0Tc3mI/jQQF6n6T3Ev8RSSLtvF/o2nUbT+rTcpl84ozX/r9nevDy9ffHE4efrUcNt57cCKopOn5q9xmUsvfI48WydcJ9u9dDKpEWk0roYx17DOXB0j0qY4bF9n2eLf/3s/PbwOb3/uP/wPiNhimS1cu2H7PtcODjJPaex512Mmb6bmw1zcHiCQuW/e9+PYNu3WUeuxNqVnXiBDOY8L7y1EMDoft7ZOMUe2EmkYHDitTm8yb/AXrzJv2+nS+gqMlfBzzDVs6k1dmcaxk0et9ziv9ejgcCAUNHkcNMCXy4M+jun4zMmj+0g1rZZlnUMO8DbhIHsxD5r7lamTjh5Kv5G2EVtXrlzJiZA+K9HDBGfryTzPhazyXlME55V4rTeC1TkmnM7Fho+c/FSfUe6Uy5khPS+dY+EPh4RLK+XR6Mvm2fyJxx4fnn/umaD0nXArS62Lv8PFSbby47zYJDLKJbeWo5fx/Sp8Lr2IpKavLNb3qai2Naz3nbLkUjh4NolfuIwhZV9gVKXOaF7b2kHrO6NTaI1jYF3jm7Z7/1Y8MOoLZ1Lwj53ioOJezlquNOGMMt1QR3mKu5yHNT6Ns9u737QchONPz7uivGxpPFWzdLBZFme3q8Ob05SmbQ3rfdOb1llvH3GZd5rCdH3DjGPHymNc5Mw33y3Ms03q7+C6wJjWaR+FTCWWIhv5nM8a+BY0UH9a/BY6zl1mDcwamDUwa2DWwKyBWQPfPhpYGjbyNH5/j5WHeLoOV48Otq9/8pOf/PyfvPed92HUfuTY2soDx/hrtcZ8f9Bzk86Jt4hRVYaWxqOnTmoExpgaIwz8oLcvcTGlCrpjci2MBW08W4QxMsdTw2IQjAwaLRPaGiDU+Rf/TomugOYR/K3gUJMWd+VEMRxlTNZPjYyuN+/6NjyMxGnnhYbmKhZb2ozOwAGgJCWrpq/GTJyIBq6c3tw4dnT7hVuPn3n+JKdtYnSvbcRB5l5P0jEiI05FImt0sUlHp5dJPUQHRJKwwT/lMq7d46eX5cnHIQ4MjSIv+5uLWziN1zb419dL3xra7lfF0tks2Yr3LgTRZ6JBlM9oE/ubaz+VkWbuXnDB33aV4y/EyL+jaQqMdWPZOvlTZwIfEWHmEMZCmxi7zhlTyaAcNVZG/WTeSIjUjr5dN2uH35dffGHYufT68O53vzt7caGyRJBgHw4HRM9o7BvVVEtHkQuaNQ/UtbqTjjKX/jXMF8swIZloFJ1+OIZkwVMwzb3ktXk7xtJglyg7DurxxReeGf7hz/7M8P1/7I8Of+SP/HFOrnyTk0XLObbLuPc8E94DLRwvk89E9khT9/AijaZHFRU1vggG7QPmEXOTqK8DnEg1E0vf4pM3HWuRyegbEG1srsUZY6SLJyJubd6KM2+Tff/qmTu7tTbcccvJ4dGnLg4rayfRl/ODpbnORSPSxv3HPB2W0x6qHMbl3LmL4uXZOmgrn3w4J438qbWbQKLPFfeIEzf/ZdyFDY5RP4DlNNXNk8NXH3+KPbu+f1i5fn3Yzp5d+4mM3LnGqbDQNELTpcvr7Fl15fIbw9NPPj2cOYUT8OzJ8HB807EB33gyp9PRsnzpbHVcnRtxiMEPWvOxKHmAclmfc6ie+5pD6tPndzE+wOkQY0kbzxpOCp63HufsQ0Ykp6crXnz5xeHzn/vcIO+333nHcBdLg3u87rjjjpxm6/tzDeei41WnWsK/fIbv0TnrS7Cf3cwpdO/8CV/e0+w8QZb8T716NhlhaeSWe1k5Pwq341VzOvyM8NLsfjUp1Q+dQHvI85yxo9wwlfscSA8gUnggz3uAvPVis/A5JVJAeYGg7enPpLa94fudnHFzgGirdv9tqj5BQ7089nsruc8K9aZEEzIJai8xyuhPujx8wVcwxXs6KOx4wdoN6Qb+gJmWg/MG6CoIY5rCel/PSsHUr3Beoz7Gfp4iizuZsat3tDyho0iEBuVQdOv8s3R+e/va+YO9nfVybmaZPQpG4DnNGviX1EBeof+SOObuswZmDcwamDUwa2DWwKyBb2cN8L3Dn6D5/aWf/9n9q2++8VU+2b+C3fCiH/p8cXNYHp/cldwROEZWL8sZHUb5yO/T8PxrfjsRNG76cg8ZjZ4uaxBqUAo7vdowahyW69JoqqU03W9qYHh/s3Fyc7tiND7bpuWmK46YGzZigGk4BneMlvxQjGHjvmQAHbE9/sH62TOnVu+5566j29gY3WgdHTuxZzHqvFduZTbSRePZ+9aBtKdl5dtxo+8Rzr7SMq/lk+QsdzNyRV7coF4abpwuv+ucjKkTxr2MvGzzin5ckpdUhqF1cUpg0oqrT+fzvpP3XZZX+5Qea0yFa511u/DRZc2jRf/G2XoVrnD1OJc12vXK7b2XfV56/gVDc4geO5/96JQvco2IhatyOV26rzRMljv3foGfZlybaZv+VD90hrG9xDHiAtBxk95v/9Ynh2ee+trw5//8f5kldk4NnSnij3wa/qNBrxNjyWfNyeazc3Emco6H0zodX55cqROgTxwUj3PC9qZj3nNtH+NfWPdGSwQZDiSX9Lkflny78f1JHMzvvOfCsME8JWB0oUuX+7azIUt/jSTzUigTjrvIpV6jW9rgLo4ReYaOV5xq5m76b/9Jklf7IlZwKbM0EWh45rnnkLTmmVGltjk3r+Mw+/znP5+91Pbpv8VS2/vuu2+4884Lw2OPPzpcfOHFwNS41Lxxm6Z2wE71K10dLyZpLMe3+qVh8tN9zU39XLburRPHLro19/m8dv3K8MgjjwzPIY/jdddddyViTFjn862caBu8wK+zvLKfC8fZN69yF73l81p6Hx1V8GJ5yptjbprWN49xjo04W47O5W9Jr56V1lvjC+LxR/ydpvQbX+cNY35zneUpn8JYzjvQdyXvOedrp+av8+7b7Tfj7/rOhfeyfyfLcAZvN9ZNcXe/7mMureaj6wtXlbp/y9gwlm/mcwrTODq337RPw5JnIvJeYXg5Q/mAI1b2D259//u/+7Z3PfDgCZ/Hm3E0D3M+a+Bb0cDyCflWes99Zg3MGpg1MGtg1sCsgVkD39Ya0DDEYscewboeHsbA/zP//r97eXf7ypNEV3yNaJNrnKKGh2xlhX20jjjpzquWP2J/uV/PBkuBrDPXUNAIyzc7hraOMhxHMeglY5SNkT3mXvu0a3x5wqHRKeO3fqIbasmSyw8x9l12yOWHfgx/jE6o5K/p/kW9DR2ddsJ4yUenbtcw1MnRBk0bDtPTC40simEKfnmWp+ZLQ1qHV9HIH/L9ozzFgtvYODYQRbaS6KDoooxbjU5OuAxPcYLBvwafLHph5uaSZ+VTpsC1kY0O1INL9Xbd1wgHRVZ6Gj7kRbLvMfZV0lGmw8AT8Fyi5bXFqXg6R+RDXtcwnrN8TyNZlfCrcyt1VGgk5qLONmVWFzo+4rxQv/CJ8KXrsJG5hHtJXdRYt77lTx2qd3no+/BMeZmcP8CCZZVTULNEcNS/fXTw6Qz7zGc/DdARjoZ7FjjhLI4FYUzidiy9arwUYpmKx5orRgtGlfDuuAgfXRkYRRdpe4GV/yoaTieGcEZPudfUNpFBv/ALPz989F/76PCh7/nQsEvkmJFo8lEOTfaxG/UVRyXPjjhtj0MJHuKMmjiQxJ/E4PQcXo1MmijoE6dP8+pIOSc6+k68HAiZuuiCe2UKPeHGuXfo6aLI/OD97xg2jzF2R5yQGfTMJ+DTR2rMCcckemAcoxgc3pkb0F4lMgxpgBz1jn5cZnkkjg1O5zTyTKcN/JvQaHBFLvTQcpg75/R87u74TpDv1eH0yZPs3bc5nGAfvbPnzhARd8tw+fKbvBd0NBNZCdO33n7b8D0f+h6Wsu4Nly5dgrdDosOYN9DuEzDlVxmcL/KaS6cg9+qmdK4CytHn2JROXfWJTkcY4ep9NjojiR7LszkOmc9xO/GffPKJ4XP/7J8Nr7/+ak4Uffd7Hhy22G9sj3faMZyGnli5Do8neWY9lbX0zjyGL+mUE455yRh4qRvEynzXYWoEnJf9+t2GAEn2z5jDt8+Vy4jVgX+s8H3Zf+jIs8kcrKjLnm+jfsAUHOoCutEfeE2Zw9SrpzqptvRoW787SlejYmwgWddJnPZv/ZuXzCV/3sOA20c++3JcOi36gif/1ozBUiW/fQtWON917aju/ubNZ8tXLNbctM5k3u2+M3xXi9OrYQI4/ljXvFk1vYciNdOreJDUSC6yGvnndcDl8Pv3qlZf84K+IupI49T73vfdZ3/11z954j/6T/5TkXIdFMruKOCcZg18Cxrw7TinWQOzBmYNzBqYNTBrYNbA21ID4we9X+i4P8pN89Uv/fOdR7/y5Wc4HewpDJFrnhKmUwKnyyFOlyP3uLJsbpvGvg4ZHTGe/qaR5tJIlwgJ52VURPer9nKm2dcr+NYryknjRyNCp8L29naira5d247xaeSVjiMtAVMbG5bbUOh78XQa5VwYMMI0juV91Wn02rfxNF7zKR7aWa1UF8t8jlYtYHmdPXsa59RmjOP9fTfKrwg6eZF3jWbrdJ5Ix0udSM9LmbyyMTd9Wsaub5h2oDX+xiGP6tSxWEf3OsoyBkSUCeNlalmk344b6zSJzVNPPk3Stq3bbbNumqcw+en2xtd9O5+A/gs6t6+Xspu8V5bHHnssRp+ROOIxOceUrWGl9/WSzrG3SuJv/TQe4TSubeskbsvSFg6/wvDwpz81fPWxrwx/9s/+2eGNS5ejPx0m+yy9M/WG8DqT27E1pSFM60jcjb9pTdszjuKBD8faze7lxav5FLf3PT+8d85YNteJ5FyUv3UEuOeu24f77r6AsC4RrKV64tABoKsDIjUXHQsF1tlCaj5DD9zhwQaNeJ15OM4838NllR7uYBSZh+M6v+2jk8Hkhv+W8Ypiy6Mz7sVN9+EE7xodY/LlOJufxeGrA+aVV17JHmTC2v9WogpdsrjJfM9zRn0/0/IWp5PvOu+Z7TqE1GOnqq+S9+FpbOxy4+0+B3gibdPBKfwOepUffTS+x776lUc5BOWl4RjLre+95x04q88gcC1Jb5wbRNidOXOm3qXcy1LPB++F69Sy6tzq+SFdYbyUxqXn7aDrtu5n3ri7j7jrHgc6c0uYr5e6jzBTOOtN5tY3XNc3vm7r8u+WT2k0vuY9eKQjq+MhFeJq/OZdnuLp+mlb3Rffra8pHdtbjm63ztRz2HpTw70VTdt6zJqPKXzfN563KjcdYRpH3RpFxnPg3DoczuJCPfnHf/AHBTN9/QGt9vl31sA3pIHaGOAbAp2BZg3MGpg1MGtg1sCsgVkD364aaAOwPuCby/HjevLhrONmb/fpJ566+L3f95GLJ7e2sPUwouOUOnAdZiygOn2ullH6se7Ja6y9jMNMnH7Ua8T3x/3CIBgNaDeKNhmpYps43FNII2dvb2W4ev3acO3qdgxc4cTjtTE6QThpE2Mb8xiDW+PRb3/bNbKbZvVrI36sNyJsxCef4V0+qTMiyuCWcpBgQBqdA3zJY740fuQ+PGGKHhklF1zgg48NjOBzZ04Nr196Iw4C+YhBjRF9RPRc+ENO9/2Z8qrsOimjD3KQSmWMrCj5yhAEDzLbV/6F172ZsAhwut+O/OhIMHpKJ92xQ/a8omzSOVQRYuJXBywhVZeEJpQzpIxcZak7e0XJcUhI00saaIk29BY9gQ3a8uw41DIxadm/MEVnI3+ls4lO1SFXMORUTJwj4Us9qX+N+mMsnbsyvPrqy8Mq+0/lNFC8ECeMViLVPNMALR3so3O6pG/0FbUWLmUveHLpwteBThsYOI7eqGJ+gUe4Ua4DHWXoiZV4gVcPiQ7b3xl+9u//veH7//AfHt73/vcPl69cj0O3nhv1XPBxzIHLORb9Raals63r1Ff4Ab88em+SD3Vk+JCn+dm2pxeGyzHcH+eFjqOCd0ykX3Olx802cXqtMV+Nwjp76tzwwQ+8b3j0V/7pqC/mDs+kmJo+yEAIEaKPktDPwMq3nB5qhfuLyStOsOzhp5xiUAadYybbR+fZqvoGp89ampzHyBenIjK5iT3+v2GFwzWNdCOaFcfPIdFkZ5gDryP30fDmpSvD1cvXcwjGhQvn46jXabi9XctxfTYOVnn+Qd1zwTFV1z7wvnYoolL1zA06DyDV3sY5WuyN78GaKzVW5eTy+Ta6sx1nmRc4IB3/J554YvjiF7+YZ+a9D75veOC97w3tq5cv5w8A7qFmJJmRi7fgzK5TTZdzInpBZ+KKmnDCJ6LIcYdB+XAeBI6y81H6JiO6MnboPnCpVabuU3AuK/aZyT6JvpR5T9Wc9/1Zc6fngH2NVJRm74kYBQJZkU2jbkda08y+Uzy2WXZOpy2zDWy+izIwpQfx2+70gzF+lNveJYt6t8Lhc34EVgBg5XMJ247R6nuYZwOwwjTm4HeOOikW9ZSdm2mK8ynNYM48F8x3Z+EpmeShk+iqXO8l64uvepf67hV59/HfmtaTY+lbyIRk0dDIdmDss4CFCR6RjD87I5xELyf3icI0ASMSwJd8pWH+mTXwTWpgdpB9kwqbwWcNzBqYNTBrYNbArIHvSA3w1eznN+lo9TqWxiunTmy9xsbiu37I17e1H9j4yGI81Ae8bbnoZr3GcZlcVS4jgG4sDdGi0GmSxEd6HFHtMLI/RtouhvrVq9eH69fqNDoNn6JnlFU50hb784QvjXyNDX7EIQ/gLuMuVYv6ZamMFWELd7X0fQwS2qSzu1PRP0I0btuzcTl1ktUWhU/8dRg5xQbG+tnhhZdfYeldGWtQWhg/0Ql9Y6igUp1YJuXQWVU3pVdM7NBdxShOm/2kgYxtBJtr3GtAG5WjXsvJJ9bSs46BdeSp+h6hMtIOxiWFU33Im5d8l9ziKp57TK3fI0xB484IndaPuan1uOSl6uxvXfMvHcsxcunX/cWho0O5THGe4SG4ePHisHft6rCFE5KTQjPf7N9zy/7RieOBPnQ6tjwa8LZZNnWeAj8uvQpf9Gt5em7dDG+7drn6e+n554avfOnzw4//7b+Bc1fH7jjuwDQec1PmCXmXp3XyI/1xiBfjmDr6Rw47ODaW0b1OjaO1ooOXueqdRyTnzAoTxhFvumngR1zWKbM69sm8cP42nFA4J5jYe2P7Cg6xAx2WltEznYZD9SMOZVLPi6ee20nKG4V2nWNxmJEfwrPLMXVE6nzyISp2fQOUXNLZh16ivSC9Dj2YioNcR+8mUYSnWIr48suv4oy8mneGkWTOQ5deuuRyyxMgwZfxhFs35GdCLPTgHl1KoR7UpToyIkvB4nznvufkYlyoi97pI16XPXtwhA4jnYnWjef9Zg7s7m0Pj375K8Obb745nDl9brj3HffFgSecjiydY2dvuSU8Odedxz1OniB5bHw36OiSB51G9uuIuD0iak3yZH3n8q2exImW8VsWv8Ev78BLh7Agy/3QAAAgAElEQVTX4K25IG2R8X5jjMQVZYz4yQJrbqo+dljWLzbdp676V5uwls07dV3mSMMvmwu+6xmU8I5+Gq94ljh9By0ji7vevMa/+LyxD1MPeuEpstrqTF46uqqGX+ZocI3/HjX+bm9Z1JhJmsJExxOZbWue7NP9woONpMJdfDUeGKBe5RQfOu5LrqJlv5QZQHPx8UyfPH361HnmwCmar1DHGsvm0B5zmjXwrWlgdpB9a3qbe80amDUwa2DWwKyBWQPfVhpYOkXegi2/vPP1rZlIxMn++sbq65yk9vretW3sVJuSjB0pc5sqo3v8YLc93+6gyId7UAmPAcDHus4q/6rvpzl/L18YDvXxj8OC/nsYmNev72DoXk0kxviBLxLK7IkUx5rGQUVCNF0dRzpojKwIn9CKEcBf4KfGiXVleJRREsT50aBg7yoML/sbJGZUi3ZE8TcadTqylJX6VZYuup9R44M8ZrfGENpL/dFwYmuTpYBrONi2o5PmRf51WiRiBvhWbWirRAi3gYNKKOo8c0z8NboMPtGpSUPOLhqOWa5GWeiW1Xph9S1oYC0jyMpZoBGcyCNo2KegMMIdT8rKVM4vdVYOMIdcfSWCBThlLl2VnryP8W6kz4hHeeJYCYUaJ/ehaz4je3AxFsjovJmebqkczhFIwe7h8CInWDIphjvO3555cYSzxfkhXJyEMLFG2ag2ekR3kpae+0dFHZa5dJDYx/FJtBh0lFsHQ3TiXBANaQ0YlyUKmwlHXe9X9uuf/NXhox/7Y8ODDz6UyMFDItdcXqkcrQfxZSkWOMUvv8EV7OP8He8jLLzQedHfJh03RruJ0+gXNIMLtcbLdvUwnbfOH2n43FmvxKLVEVUya+o4qPyPs+ccy4PxtQ1XdLaylx2Uas6jk/R3zkZxjO/hriTDo2OmojJfkfOIORIZbHfgnCc8N2p/oQfm36rzJM5zMKCT8MJbJm8LIttuOXtuYHXlsEpo3LEs+6uxwh083HJma9g6sTFc394dLl+9Frw6hBwel2NKx7HLOEKjHagZPuaMY28qp1g9z84Knd8VLercLhikD15UtNCDMrmk0rFc6Jz2PXTnPLXv1554cnj00a9kvO6///7hrnvvYZnl8eHqm1dSt7ZxIkugT7K/2qmtk+FxJIkO0eN4IquqEd8BkXu+D5NwzLrk/GCkJw/eW+f8cMn7LUTgefAATDJ3fK5qrrhfWbxDIOIJwSmK3JmPVDDAjrv4BGsd9DyWts6a6Gihn3qqUPdCr3o9875E4fb1cs6Zd/Id1in1LTwvv4zd+C7uZ8X5VdFWhW+CKuPguyvPFLl8J5rM6Qd7zi5204wO/IdM51j/0UEehJef9Kfss1rvEOdA3Oxx8jq29kWQnAJrbvLEV09szYmdoxzqaGxeyC2d1gNPAONM/+hT2s694l2cVfa5lVfASs2Zd05f+4rLOTgmXsm13Jrx29zd27kDx+kdtF3nQj3FK/cl1NhpzmYNfDMamB1k34y2ZthZA7MGZg3MGpg1MGvgO1ED/dXsdz8fzof7H/zgB1/b29t5lW/v6zo8Kh36/Y/PpT7KNaD8OI8B1UaCuZeGNHk7WAITJGV0StA6I0h2dnaH6ziSjBrTSSZejUxzk4ZtO0DKAMYIwXBq2oVbjJUs+9/NSXxpC90lfBsrDR8jYtkcOXSaHWAdQznOmsaevuC1TztatPncg+3UyRPDFZZ+SVPaXjoLLQvvEjmjWNqpI33bytFTutXwMToFpaaPESQaneISh0vOhOl+jSP4gfEQBXUsTnXIcAWXZY3cOMmsItlHvekwgCoVApcilPPmJE2QLMap5TKXJ/tE5+aMZ4xc2tJvgqzL0u/UdS2bZXEdxwHy+Fe/GrB77rknPEun+RNHX2VIh8WJnLQzN1fRSemw5lfTbjzhG5rlJHQ6K1PJIHH5Uh4s8OHliy8On/70w8Nf+sv/PcuCr1vFmNZcE2/RKaO35y/okpSraTff1TI6bBzsMTWu6MJq1CW/HqzAjMi8hFigc+gAz6ljmUMxkNlUDk3GAMPdJG/OP9c6H7HMzyWrp0+eGi5fgy9wF0+jcw3nhFE6WV69gnNMw5604smPeo6YO3lXHKG1sW8BxB3HLXz6XtDJYfQWjij9aEc4E41acryghEN3lJnnw+WGiqQz/vghc51DBFz+B8ORy43tV7eIKDuBF435mvnCW0y+ve+kY1odLeaK7zDILMpjW49Bzz/Ldd/zXBnBjTPE53Jvt2joKFOP6l1ntUtW33jjjZy0afSYS0XPX7idDfjP4DTfzembcYqdOcd+ZGfjJJNXDzU5vsopluAwlSNq+b6VhuNttNgbHEIgbpPzypM9lVkHmn9oMLpSGscP17IEWb6nr0WdP8ofpyu5Y5AxCsbSTevBKu+X+qjyCJr6KUzqx2F0jnUKDxTMdUb5vw46n7NOefacKySdmKs6u3lXST/8ktuxeBOPaXxeqA+PmYsgH5OwdgtubkI/FehA2vxfyxrHOT/OwZZZZ5l9vEyhQf9EtZLHkWauSKpypFt3SydZ4yveF0C5mdY1Hf8YYX1fUu97O3nvmKsXZIuQuvLKkTicQGN34TBlo8ZjL/Ev9xXhwV3KhdUQnn9mDXyTGpgdZN+kwmbwWQOzBmYNzBqYNTBr4DtAA/0Ff+MnsrZCWl588cXth95/9DonL17TSM1eNjE8R6MFMLv2h7ydNBI0dvKxPhoSHY0ksB/nttnHS7tpH0PTSJttnWPsOXYd43GZdISVceByo+MYwzp5ykAofBpGlUbjKX+xr7oYD5SlKf2mHXgMIPnXDpVVDae0l9lGZSmoeWYLozgMNIo1gvxTfkWZcBvDf+RCZwVyupzxFBv1x2Bf2cMRYCe7jfJrlgG3g9Ml8rSxOtKXZb0HOtCk5x5FyXWQwfA+cqWfBjMw4QuWNSRDZ9S1MOrMZXPyZF+qqq8iRpbRqByNwvTHZHUm2N/UY2ZZPekkDS7aEiE4wlQbyhJGxZJW0O3NeNwXy34yE9wBZKzZK01YsI90qq8wSThNXEpnuu02lgPiGFhBLp1VXjou4ohTz42bvv5XxjFOGceauhrvkk0+3APPOpMOGfGoz8iaWp2HrV/kY+yMevrkr31ieM973jO8+4EHhh0OldAhqQyRg6WJu0SdlXNS2UTEcwIaZTombJ6lnschVNQA9vkRLrqitvZMKudA9OaYgUu+OTECO1ie6afOqdPR2ZFx1it79KMzCpKIXLpZwfnHnNoi8lGdHhIdBrrA6uzLuMqVz0Xsa+hB64jxMgoxKR0o6zcUOe1dL22F1znGTarrmTOCDL7QY6LOHCfGMDipO8FSSh77RdKDL3w7lbOsjrKOwMwZ988iBbcnclJv4hHhvpbxGlClCEKWMw6kjgKZY+Ec0nln33JQ6bZjPnH5vnI+OC4urXRZJYfYMr4+18eIKORZR/Yrl68ROfbo8PjjjxNJupm5eu7cLew5Vo6zM+yhduHCheh6i3YP1MhBGji8dSfKXT3L3IPfS/42iKLz4JLr167lYAKdcB7C8forr8ZZJh9Gjl169bVhA5zXgDOKzFTRU/V8tF7MoZT5rrO953c/b5l7zKOeN+b2iX6pl69MCcee1Hjt1/d6IoXv9uB2OvBf8NBg5G3m2IjfNvkaOzHXGnf1iVMWGoc49cQXnEwOn6eUxZ/xW2ApJ5azRFZpE04K8l+zh2elaRblwAY3MObOP8e/HGYlk/U6LRfypi86gzffMyb/rZjKR421mUfdz1xuxRcWIea8pesiya9M6ej23xYdaN7LE4kpw1J/BSLhyF7fPzy6Y23j5B302aDmStG9SchAzz+zBr5xDdRb9huHnyFnDcwamDUwa2DWwKyBWQPfcRrIR3p/V2MgP/yp3zIy5tLR/v4bLs3xQ50MmxtTXcPDD3IMY4223hRZ55gpBgV5ffCnKj+Wu03DyCgIN+LXmLzKpuYaftb3ZSf7aND31XXW933jNA9NDDeNEcv2a7hp3vdNq3mzj3VTXLZ5YTInt2/BLWXtfumrUwKT+iR7JB3HoLVOY6b7Cdvw4jWZNy86Q+S/eNc6KqeGfXQMqDfxeVn2sk0c5mU4La0q8YpPg9u870Obuu5rudqWPIW5yY+wXjfDTcvedwoNCuYtn/2n98JO4ZqP1lnzHz7RxTPPPGWH4fY774jsTbv5snwzDXH21eMojMncS30L0+XQpex46HBqh599bHMctq+9OXzhi48MH//4xyv60WEuYzUwRGEGn3h7DnvfSTwm876XfpULqnmq0nLONU5zZW7+j7XDEE/QtK94O6lby45U9OfsBo8b/u8Q/XQMZ4mpxoCxi9Fdc0d4vQouAVykUY543PS6kXw3JI3yhj794iSmq0vBcuqjHgBhjCyDI94qcSgSWkoU1Bn4tLn0F4cBFZZN5j3bnN9dL4ut7zjXcWD4JljXCcQ461Q272S/1nvjsOy9BzPUM1W6359EjiFFYBwvnWY6zIwq6+gxHVSeTHnPffcGrpc/6hw7zSmcOnl1jDX9jAU0jfpTcHloPoTR0WpZvG+89nqcYzpnnnnqafbA+zJ8HmU/Nt/J8hSN0q/x6yTM+CF45gu6PYZTzT9EmMR9c7LOPt3WuThzjV28d+53u7lRYjeUe55MiDSehuumTDkKwYuedTwLU+V6ZlLWa6WjeEyNz/xmnN0maN/Ldt/zDxuF5btTOHE0nul94zfv1PfBgBe24OsZ8149tv47n+IOHh+c0fFX5XJKNu7mwXLPYe+58JHXQykMy783ye9kbO9EPzjIFnL5yCyZbubnfNbAN6iBfud+g+Az2KyBWQOzBmYNzBqYNTBr4DtAAxo1o2Ejt5gAZlgUfEYTrfR//C//8/Cjf+JHrj7/wrOX+PY+WMOg5C/SqxiKBASV8eVH+KHryUYniwgWCUOpjGudaC75KCPDun02EjdqbIcN8K9cuYKxdx2jfC8Gpiz413A//L3cG8xL8/YYBrWGr7g0iEajoKJH4MWym5bnomzK3mfcyqtJfgGJPdU2lf1M5lOjpeUMXmzpQz2E0C768EhUm0bcjUZgOzrYz4klTpvrG1nypHGn8apLwksckQW2FMcT+jzhkgZ4LF6lq+ymMsC9KefJ7nWcZBjiOmkSxUJ/o/xMynqAjo3ikT9l0iFgdIL9dfi0rOZ9n860V508lvFv2VS6sc6ldgW3GA/aG07YzA3pj3DhZTSOlUU77sBTPZk+izYKGvQ6X8XVzgDxqTujjDhglaVlrw0r7D11++232xTdGBIkTnn0KhmqPOVLp263y1v0AXzubTPSYwzZKHlLlu6DFkLTvZ72cX598UufGz70oQ8OH/jA98B5OZVKzOUzUnOm9KxM8mOUR2xx0OlG0LliCh+5I1pp1F/X2a/A0J038B0Yhqdl1Dnm/dq6z0s5zezvsr/Qde4jX41o9eu+KziPtnkmd9G/uMMPOnW8kqTvFPJESOY+iKreX9poUYDo1Lx1ykBnjAVrnepudrP+Cg1ijjM/dZwlcovoLTgeCIUa7rn7QqI8paUDXl715SSyknvZzEEBIs/Y6Ezw2Sp5DShrNjOfYc/nzQhGRqjkAW90BD7xe99XVo4GL6eFUkjUGGNvKqcZSyvRj9GHlrd5Lj1E4pFHHhmeeuqpRHPdc9894F0drvEHAN93W1tbmbvnbjlTDi7GTB23s0PatSdiOTHlyctTSn1m9D/qhEsUKWNlX5dUnjx5mghGTq1EtydOnOQgg63wGV1Qtwd/ptCCH99/Osd6TKyXjqmW6PnuQYFezolctI/3RvqVDhx254m4x3u4yCzTX+NFatzSaf1a732ckOBoPPuHROI54nTViSqMqfoWXctd33kizWA7FOnTurO96dvPOZE/8ow4un/8S3FsCcVzxtzwMgLMq8URfoqz6dgr+hwdbUv4wqfu7Oe/cR5CseRJjtUZChznoD16TPw3wUv45tV2qkgL/XJDvChjG74PDjZ4Fu5g2lzgRYsXVljRZ5DHUtXNv7MGvhkN+FaY06yBWQOzBmYNzBqYNTBr4O2vAb7dEVJTh2Vrw/DSC89e+/Snf/tlPvhf8aMck/M439aYx3ys851ehkMZLhoyXtME/LSYj32NOzc6v3ZtO1Fju7s6dmqTa2mEzmjcaujqUGhnWRtyft97Sc+lVd5329R4kLhtb5W/VZ3GyJSXdORnylf3s074MtimhkvxU4bN0SI6RMNI3B3t1fcLehqhylQWT/iW9yxtNdc4g579D3BgmrqvuZd7D/W9OgvfDFTxUtEG+CFIZQg3rdSAW3rRJeN2HOu5282tr/ISzn7WTce9cXSfKW7vbTcVrsqrrhwEN/fvcTVXjt0dlpa96bKykywdu90oicwP+wnT8MJ2avkbd9d3WYeJ96bmSzyRTfnGMdGRp34tC379+tXh4YcfHn7wB39w2MbhW/1rXmroO1Y+S0YILfYeG3E1PXlrXq1r/nWASUcDu/lsflKG5+YrhPmxPrJq/TPfCh/La9cIHiGJWwfkIvkEj3RWWUaNV2b42gsvDldwsuCPDK6mIS49VYFvBCOqOHbBrWGeRB74eD/1gMos3cc5qbPOvbqS0Oci4aDTMaOzM84zGs6cPsV8b4hxTLsv1eq503KvxKoJD2Oj91NZLHupk4br9sUY+J4bx8cIOu/r4AXpVpvovddx5fOnw1oH2eOPPZp9984QAedJlaeIIhOv7efPny8HJvpwXhjhts6BBDo1i59aCipf7TSD+OLZdkmlOHXACy/9u+66Z3jooYcSkXbfffflRe5Sy42tE7nPvACf8zeJSW8/L2kU3dJJ66Pz6jB2A4cOs26Ls7znAbik81YpOlo8OzUW1oln2qd5Eof3/luTHLbl3X8TLE+T/att5N9ZDt6+hO/7zru/ZZ6cLt6A237dtwEW+rPXhEa3dx/L3e699Z0a59Jxu6Rvn8bR98rXfaa5Y/ZW4waPKITFlwcH6zvXty8wH+58/wc/GG/piHtJsJma81kD34QGZgfZN6GsGXTWwKyBWQOzBmYNzBr4NtXAjXbAv8hkfb/7yzc0hjOOh2F/d3drfeOlg939lzCidjhtDixZY5m/pxuK0R/v44d3DJXUAantqgG7vI7iHHMfnt0dIsiIBkr0E9jcdF9bpSOddFp4EqFLf7ADaJO1MhRk3rL1bSBIf5o0LmwzNW9VgB9tOA1evQDeaghRR4/kae/6xqscwowGTAx54BOlo0MAVF6Fq2krk6cZIucYdWK7RlYiosBnuXkQpxuge5nUoxE2yqERa1mDkX1l6L8Hzt04iHQSpc328QIiOIwWG2/S94BNwK3yMhKn5Wk9WvYyubdNRes4hjrG6BNjsugEbnRWRK6Y4oXTPbykbS42pczV8hItp2NFPuW5x8p7k0OnjDpIdSKYXHZ27fqbww6OqVtvI7Jo7QQRMzgMGUdpeTX/4pMno0S8b7wlG20iBF59ejl2cupcLRaca8WbfZme8OI4OA+QH96+8IUvDMc31oe7WT63vcvhEvZH2KYtCZ0U7u2U+QE95xAjigOIOQfOzDU6taO3HABGORbf8utTJ5f6n8pxWU7KjkZRzjyz8BuJsI8jNzLJuziMvmzdRGIIZ8zoC8RwHAeNe+U/8oXHhu0DRplTHpXFPspjbqrc58S5uZwrtlmX5wKdi9toPWFATyMj7TPAfMm4UJ+c8Y0iAlIyL/SHw+jMmVM4j+wOLvryG30kwkgeSKgllxFW3qtLNEw+8iEQqeXvuSB9o6BWGIhuazjbvEx4G1A1zxhXLUWs59Bn0mfwYHSMXb58ZXjuueeGL37xi+yT9/Jw2/lbhu/93g8Od955YVjnVE2XkN91x+3DHbezd55LPRnQ48ynjbX1YYujOl0q6bvBd0VOwuTevcnWDYMjhV9kFubcrWeHu+6+e9jAUexYPfje9w7f9e53D/e98/7hxKmTwzvf/V3D6XNn897oJfLuUecc90qUKnpayANe8euYLa0WPeetfNY7aXym6KfqveK451XjHz4SfcX7ymFv/TmHfL6E7Xem9+XY9Llk7Mb3Xes7soKHtwLt9a7xPdE4bU/0F4S6T89RJLIZitBFFvlX3tRRXuKouWa557YwfY+INanIwgMYldXUNK1vutaHFnMw9zwDKkI+885knPPMFyvQAV4uabefHIdmeltEdl/hzs2WCV5NU5573o58uwWCIGr7QHf44dGxc3fd845b//Enfm3rz/y5PyfRG9OkPLm9EWYuzRq4SQM1y2+qnIuzBmYNzBqYNTBrYNbArIG3oQb8Ai8rwOzoYJvT117AiHweo8xj4sfEArF84S8/qf1ob8NzmlvvZXSFy3+MwIgBODp1ut1cnObZjJ+oCo036/zm1xj1vq6lodd9zE1d9l4+LI9Gg1Up5+ame2GahymO5m+KP0ZR2SpBJR3hYsCrNu51Ogi3jnUfI5QlN41D+OYp/eRFJ4pG8yiniBu+eZj2UYcayuJq+qE7ypzli/AhjPU6mtRjHJDcTD9wG6/0mmbZWDcaoMLZLr42Oqd8dpt1puZ7iXNZ37issV0+vUxwXDSg17LpOAKMqMM38dvuDGfO3cqqPPduqqW46q1Ty2NZ3JY18m/mY9quIe9lEl7ehfcSt2WTPO5C/9q1K8M//ae/PnzsYx/DmWFky43zT+NWw3aKQx46df2inxoFh46DqW6aJ/t1hJSOjjiMqNO4LgN7nHeM/zQVzuVktSwfU/mM6DrGRvHPv3pp+MJXnsCQP56lhD1+2TRfpDgohU1CRzBcTjTvTeEfWurKa6xfNWxx1J9OtOjXsdahRx/7mVJPLl3vGfyFc1QZM0dcejfOceeEKTjy2qr52rKlkZ+Ww9y01G/R7fpuA0vmoGWdIuKXpim40YE4us56D9HY4d128aUXhq89+ViiwnSM3XHn7VlG6fPqiZJ33HFHnsVsyM+7QTwbOFl9Pk39DJRMNU7OPy/rvKIbYI0kcw8zry0i7YwCFK/1LuM8eeoEz0g51qUvvzr7fE+JIzjH8eyyPEz1IT3L0zphrFdPOnBycufIm/UmaU37Nc+2NUznwnnfedcL23WNa4q363TMTfsYyWjZKzyOTvyua9hy+hdc6pClaeZm8nOUkMob+WmZGq/PauO2re+bT9F1feQYy/azbJrCpmJSZ9s0id+6zrsdGrwqWMSZcVs5tn9weI5n8OQP/fCPpHvzNcU1388a+GY0UG+rb6bHDDtrYNbArIFZA7MGZg3MGvh208CN39a/G3d8cdtMh431bb60X2Cfmhf4yN5Jbf3V3hVH2YsMMyBRMJhQwenePhoo9cHPkiL27fFDPcZtnCC1THD5Ya9hQG9parjR132IVo3UGQ0O8bkcJdFIRtZgGMSUMdINoDge6BucwMEa92XYWmdqo6DpWtdt5m2gWG8yWKB6Vt8VKqSrHeOeRyvuMWM/aY3yyrtOjBg/RJusxTnWhm21HccJVgrWWDXKpT41acXRoa6Ek7IKyUCEd6NcFvup4VyEDNEBmLtZp+MJn2X8HiOaJBFVYtcHwUl+R4xBTrEkEiv7azFG0vDSYCt6Sk0ajUk2mqp9eqxDXoD8H6zLPofOBYfPduqRNP2DN3V2cz7Yv5whjlcbdOY9Ln2f+SM2VeB8AK+49QIZIfTCs88NbOY03HrreeYIDoa1fXLkos0rfDJITJ/grtVGLiODFvgOZFXdkLvxfk4/jN5RFqn5cSwDmlpYCRtE7+Ho1dn75S9/cTh95uTwfd/3fYObth9f7Sg3NcS8MNqIyJ84yaAr3sznBVaxl+OlaapP+bJekWsOI5N91WMhiHOyuJUp4cwLJmPA/YHOI/Xu+JCcl03H58ku6sNlfesnt4aD4+vDk88+Prx2+epwnKitcnrQ3UhSUp6PkQ91ecgBAIlwCW6QxcCHR8dAuHTix3mKc2Z1cyPPzeroCEqk3MizD/Mx9uoz4ibvExxqHT0jGlN4B2/GOM41nzxSPJHU4+hZzDWqdbI6ZvYLzryX1Kujw3/wZX/b1fMYTMqUKzw6XXSO+SzRafH+6tMtow+jf4yYAu4qc9KN+Y0eu4YT9/wd54cH3vueOPg8gOT6lavDO9/5rmENB1Y5sTYzn5XiOFFi8i4fRpbVMmgjFj09GEng1XdO9p1DTqOSnF/uU7ZxYn3Y5HLzfyMtjcz1ubFeOnnvEhq4spYRQX86e8dJgWTRJ7jtk2d71Ikjgdgk3yM6NXsMxmr0pK6c1HFNe8wvKbhBx4yPbtuxJx6fxZKlcNlD+sputJf3Xc4ef8ybNWSkMbgcq3o+LKsv+oHEsXC6O87izHjKvHzQp3UbruDZujTyO0oTHEU7lemjbD7bIvW9BTkSfXWkWXBcigjvWauKZiLXRlD5qiRNHKn90MCDfFibPfSMmAtfPgaOxMhh6ni/qGv+zSlYbumYf2cyNvUHADTMWGV2hzV540xL3n3rJyG7tXXiFMTEA6OrUaACLFLd0p6kJuc0a+CtNdCz5K1b59pZA7MGZg3MGpg1MGtg1sDbRwN+Iy++jDFutu++++4XMK5fpH7HD3I/3blih2iSlJFCDd/cMRDyya9CWC5EnX000qYRT7Z2P+9NlpcGUhnzGohlzGgQlEGhEaTRoYEkvMaTKcbCyIO4pv0se5m6vuFTyU+3T8vCmKZtZacs8S3g4U/oxm9uP/M64GBp/NlH3qfyWde6ilE88tz41jgNU4NXg9OoNOuFazlcxum9ByCoa2l3m7iF13nSBqvt3d+2pmO9VyfrLbupvMmyeE09XrZM+6dPIOpnis972wMz0un2brNX9qmivdsc8w2Wqb368isSG05uebohlDEs5aPxNW5x2Ld5FdTytE5dNNwR3pRDDVBgxGGyb+Od6mp3d3v4xV/8xeGjH/1oDOjGk072I6KseVroW1YncjfezkulZXbAAnwIP35I72gAACAASURBVDprKDjvTepBHmMsYwbjio6TzzZplkNnab4ElrbI5bNiX2GRXfjMQe736fI5osfWt07jGx33rwNW/uhUufwDq/NssYdYZCo9ilfskhA/nayiUJvQeysfmd86uWgPf6NzqyMHXXYtb0zkYYvINh8s3zvFi910Ko1LRgGLMx28rfO8G0rM6C2yNy8yQRKHV49x1daYh4+R9YYRbkSZzfHDd5xK9FQf0P/a177Gvo3PZ57ec9/diRiTz9dee439wm4ZbrnlluwbZoRX9a+9x1xebnlvD52Mqfmz2Pc+9zrB3Fcse5fh3Dx16tSwRWSaUWRGqJ0+ewoaZ1Lv3KsI1uVYZ9x0so36SK6uRzrm8tLtljMW3pDCd93m/uu12b/Ho/vZ9+b+I6oFPdvVtU7o4GDei0dZGl/nUx4bT+PvNsuOp2Uvy17d3rx1e+PpZ8+yPrLMWfqZmoZ8dOo6eX+rNKXX7fbR4Xcz7Sl/N+ObwgrX7x4whS/L3d9cvona3lrb2Dx3+5138jAlySRKGEtzNmvgm9TAHEH2TSpsBp81MGtg1sCsgVkDswa+YzWgBeCVT+fNtfUdHBIX33n/ey7yNb17hEFgJAqOryN2AI61oIHuR3sibkYjRBtBc1JD1y/xNm6FwzxJtIAf7/UhL85DoiF6jySXU2IQaXxg0Lvvk4ZIoiomf0HHbAubK0azQFAHgvikJp1O4W1iyFhv3RSmYav/sn0K123CapCvEmHVxosyViSSxhj94UMONNTdgPsgS9P8pFR+OdXoK6eBUTziFpe5zi3lNUqnjR86xmG0StTOJnsVue/RcYxj9oTLktU2JsWxf8RpmESMqbfjR8eD7xgReZ2E8QQ1/xN/ORrloSEqV/bwBVzuoaWMdM8M6RPY7N9RI6WjMhq997Kv8lTZKMDCWwZoyVzt5RQpHOpQnS5xJTIKnV8mwsmxP3nqTOaW+DUyZd/7ThrFphVll5cKPSESA/r8lz2lEMYIIJ0Y+yyRUzeOjQg5q5U5LWL0KFodaArP9YlPfGLYYQ+yD3zoe2usdGRFD8BIFxnlXbl6nztH3WfEJ6IdOpKCw2RGA05THHrgEiQ6gRfls+wv8SaRoySPiLSgL56dkr3mZ+tEJ23rVqM5J8My/sp+SCTeq1cOh8efeWFww68Y7fIOT85PhBv7lmxRJfqRFkxBltwLvOozzk1zadouZ8Gno5VChOB5AG9g4TtzAMfikc/+aOSvsn9b5jHBeYd74IekMvhuCJoRd+uYVpDXnAtN6cjySNu+XurEABqTUX7ele+QO8bbuSmMsLvskxgdOk/gzTmQPejg3eicPSK53rh8eXj+uWeGz/zOb+f+ofc9ONx//7sSFffsM8/n5Mr3PPi+4RadWDjHTEadbSJnHF3wt8Nzr9zt+PNNIl3fi3nu0Lfvkg34k4f1dZZU0g/p4gRxvzWT+rbdMS6nTjnSN4xSA6fvFWk4rP1+EX+6I69jo9wqm+rx3mGWrvXqxbL3RkTVCQoZV1vptNCx4wSwfDi7dWjLsjCRjZxXlb1GXnES+m8G/Muj/IlXOdMH/Stx4xeOxYS0E2nHOBjpJi4T3NYtNE35t8sbZSKz35RX57SngtZ7HABwOfelEbkVmmSfujFeC9rohUpbqp7f0l/BCpM+9O/65r87dNlcetO0oDet5F71599IogNHERO9ecQYpQ8vr7QDB94N9ki8bePE5i0w/AI9Rk+sPKd3hLOf/3aZbuQiVfPPrIGFBnwO5zRrYNbArIFZA7MGZg3MGvj/gwbq61gvDnYo0QlH3/XOd728s7P3EsJfibHADR/c2BujscgH9fQjXr/Z9EPfe1PXdd6GgOUy9AJVRhG420GUj3Y+3GMsUd/GUpCOeIVpfM1L5+L3mibL03bvuzzFL1xkjpFUJsNbwcaAHQ2bxmPfMlDL6dX0mxedWh3pdXOb/YwmEcYrBmaW7JVx6/5Cbt6tce3VfPZhAEUbY3Pc500cJmWzzbz12fy23M1fy9m57Z26znLgMSQb7xSmlulVW4+PcF7ikIfGZS5Mt6mbxm+byQi6LLFkeho541xrHL10s8vpMP7Yv+ULjdH5IKypacZRYJn2hl8ZbUkdbOrx6tWrwz/+5X80/OiP/mh0L1zrRjymqUy2xSFB3nSEafw6W6b1tpmycXwtXku5jWAdKzqpu48OqcCPOlI+6dvuZVrClh6lrexe8raxuTY8gXPslTeuac7DHGPBHR3TP/ovT0XVi5MrcgNeJjY16tO5AE/1CqGOMgObsRVPz4MV5i+MAsu8gk47hnsOiFO+5XFkI7yEZu74sf/Ekm/ckTt6Kv4Fb7zeRz/ktrqcLQ5jiDS0tIW3reihLw4xiEPQfvEQGuC2P1zfvja88fprw+c+98jwysUXh7PnTg/3coqke4Jdu0Ybyy7vvPNOluN62ADOxxHnwgGEyjx8Qp5bNu/lJXLII2V57qvHzdw+iRLjPeDyVctex9iPbI29zYw89aAIk/1tM7evDhTvOzU9y33f7a0/875vmO7fuTRMwuXdNenTMNP2hlGfPQ/Uj8srs9wefOYm+ZleTLDUd1sXGmZa37LIt/fN//S+6momyJePf8OZ9719Ws6m2W1d7rzrm37n3W7euM3VW8N4j9QLmbtPt6/gNNXhnvLYF75W4H3lwD+E8PxxvwmW24E5v7J23CNt8aPGw+ngLydAI5/zWQO/hwbmCLLfQ0Fz86yBWQOzBmYNzBqYNfC20wBf3UerF198af/zn//i7oe/7yOv8hV+WSnHD3P+0Lx0TuQTnu/tRBJRGGHyV25MsNEI1QjwY11oatkby/2NNAA0NOKcGI0fT08Uh/uuGDmmvSW9Nkhsa4NC/KGX730Nm/re17ix3st+ZWgoQfFn/07eBwcV03vrNJZFvaojQv4Dg61M5Mm+S6IQp8zZMmQj28hf09SZs0OE0n54KsNRx4B8aRA2bfnR4XFwUKd7Dvi19FTGwcIauBjV7Fm2TkjTETbvyg6y4UTRcXOMPbDCI5tsuVeZ0XvDLhERq+sY0LVHlwb+EREHGseHo5OlnEIKWTptXhZ6wMhKJBHt4Y+xQKt4B0pXDGRpHB3pOIg/ZNSnPhV1I87oknq1rtzZ/ws+dMXoIAjukQfvwyNzw2hCk5EaOqdeeIEoJ4xnnYTqAwgU7zAYOYXhD6y0DuFFjt0rLrQFSkU5pMRptJAcmnJHv0UkZGqdq+Igwoyx0wH5q5/45eHee+8e/o0f+eFEBrn3mHPNsfbSsRUc6lo9wJmjlH2J1AP4lD030RMcRC/qBl40akOTH24Wess8s8E6nUY6ybgX2AeEJB5vbVMPFa3HuNpGfaL2xuWfjoHX5hYHHWwNw6d+5zMOaaKinPM6BpzvLj2VJ5NjYjRkEm2Z38gEoAO0gLNd3Brn6SlMZKWPTEd4M/QBziTbgRZnUePJZnyd22trG8PetnTECxQAOcUwNaKmAvlCk9vogfmSaJroo+Zg4Ohjrl6N7pFWItDAG13T7wAd5ZCL8Ake6vYJdbp+/ToHRJRj27nn6ZAHHNjwxqXXcJK9GkfUO9/5zix1vHZ1e3iZ5cB33XvP8L73vW84xf5P8sdPck+uPOZzrOMV3OGZNnlQBx5UAmfcl951BCbajgphwity1J5i8AGAp776PhBXotzsnISk8Or4d5KX4FEXo85sK0dz1ElBDVWf5qv7Oce817kYuUbEwnVSjn42Qos29R3+mMMVkVay+2+HPps47nwvwJdJ3MLzE36tK176/W4NyQmeLuPz7fM/8lLd4QsdOJ1N0i6eqmx9+BrnpjFvmd8BZl7CW8tglffCd15YRhYmOgAgeNRiwzaeyDV2tM70Vm3CORI+j7qehXETUJP6TaQr977/j1ZaL2hTwUl4w/TM3kb5Norr6GrH8VNDWXJLZd4jAs9p1sA3oIHZQfYNKGkGmTUwa2DWwKyBWQOzBt5WGvDrnw/sg+Hxxx8ffv+/8v2XcORcOo6jZTSM/PjOJv39EY5FFoPhOM4EP+D9aP/dnFTdrw0CtVf3GDEYcnGOYRxpcjSMfbyfpsZjXbf/bjA3t9mv8Xtvajx9Lz9loGDA4bETXgdT4RqNJOo0SuXX/ovIB2RwTyCjarZxsGh4b2/vcngBSyHBoRHf9Mr4LEcYTdGfbTrRTBpsayyH0zgPDXBfX92NUelm0jHo1srgHlY57Q9D8xhOPJepaXjax9zUMuvXMOm4aD6q5sbfbBBuFXAm+8tvjHu9mDqgSPJgm7huTl0fGPoWjHhqrggvjO3NpzQiF206AV599VVuDhNBFlidUyOhm/tazhIs8n1walO2jPoPqSaVA2CVeYtbMXOv6C3lSLAFjrZXX355+KVf+qXhL/xX/wVjuL003sGigSk954dJ6eXdO/tLS2dGPxPyMdXR9D4RiSIhNVw5lnCWMJaVytHCwAFTcrrJt/DywU3y8VYjOeVj49yRP6OijuF8urw7cHrlYxx4cHLYo2vkd/zsrCROEvRlfU5FZDq6Gb84qx2eWOamEuKiHGkVzz4vzFfbSfKWgyicJ0ZlkVr2fZ0W8k2dEVB7wFzdvo7eNqLLQ51YOEJ0qAqTRF0cYRTU7TGWJJoaZ98HPrR1dthe7yv99a2v+O6R18hEl4eK75VXXh2+8tVHhyeffDIO0egGPl3uqJP2/vvvx3F2dbj9zjuGTQ47OE4kl0693csVDfXggw8OZ8+eHTYSuCPd2nw/zyOOOJcUxgmoUwj+pGmKrnuoKTt3PSCilx3bLrx5LWXnOUCmXm5qvZeuFZPjokNO56pO55qb4qjny/JUZ9EJveTXZFs/k95X/5rjwnbf5smylzx0msIoZ8HUe7Rxe8iIOOCqu1X5LfgTdUffNb3uZHkqU2iHJyEY39FZaL28tDzdv3Pf0SbhSifjfPG5mKRpe99nDMZ+1k3TzeVus97LvvLUurUc+ouJXz100qotJ4j97IM8iAc0elSvvH82aLudaOML1HC/dznPtF3HZN9OzJK+nfNZA2+pgdlB9pZqmStnDcwamDUwa2DWwKyBt7UG+F7W6P8f/6e/Mnzp0a9u/4X/5r+9gtNnFwN2HZtulQ3N8xXdBlDZ7bUE0KgIIxY0PPJRj6LKSeBHuIZpRdyovxja5BqAcSrxcd59/GjvZUBd17l9YwBh1dbH/fID33LDTe+tK9gycvr+ZmMkeEeDwVMm5de+LmURFpNDzuU6fDeewFCnaWedF/ZKIkvcJ+fUqdO00BMDVQeZhvHONaLFyK8RnSLuQ5VLp821zdA9xKFmCl2MHfchs/3Ysc30RwvD9soOVKtfG3tu1i/9QxwNwmeDb4x+9RznXg3fYvmWMNIwte6iL/jXKO+IFB2fwrV8GmAZZ/pbl1MMxRFM8q0uLJQc2RcnbUvrX5joDhydSncY8lRkGSk8bL+2nSgyhE9koXuwuaxMmY5yit5oUIIQLnGOla7CF44B+VRfcpeIGnke9WQkxSGOopXVWu6GYuIMytIuBDBy6Cd/8ieH9zz4wPDh3/f7weUcK51NeWUERxFGWcSrXqSZpXQl60LXPg/8h1pr7y+cL+qqInl8Fkqm1h8+EHhsHDj0xKxTjm7qXHj5yQma1GW8EXsRsYcedEiqak//PL51fPjsZ54Y3rxOuOJp9/wi2MQ5N4ba6HyKykap2HtQIugParlA5AB7OTdkRBVouDNO/ChNesdhJpPM/+xP1nAKTwo8Aq6y/PKQva1WOJThtUtv4HQ6x2mt6DpRQs59nJk8M8pZZJWnnm3rgmtUv3ru+SwwoxonkhFE8tptOnp5yhMpePXqtfxh4JlnnoHW6nDixAaOsPuGM2fY/P70Vub/yy9dHD772UeGv/uTP5VN8x94z3uHWzhZ9dKlS9knz4McHnjggeH2W2/Ls7fB86yDV34qOkyHnnuc1fJn69sR7vLyer0ylkQEqee8UxlM3cE67PV7KbNcK7POMfGxkVbkd0+u6AI5fbZXj5vrHHMvtThNKAsKPvB4X1FV6Z6+qtL5k2fTfwyA1cHWz2rrunrUb7/zlScXTsDoGD2a4uDLePtvQLXJU3iECZ3Dpp7/dV//lvS9uVNH/FMevPc96IOgQ7DahZYuP6Ua+nDL/Ky+NEBXWHnIH0LsAEy9LyzUHGpa5cBezh0hOvme7DllXUd3wUFwGtEqnoYZH7PMjcZhm/z7rPuOUz/+m5PIVIVTDnDUO9vnQm1YVXipZ5j6vZHxW9/bPbj9yuVrt8OfSyyTfD0yrHQbFUNtULeiRrg5mzVwswZmB9nNGpnLswZmDcwamDUwa2DWwNtdA/UJzsc+IU/DL/7CP9z9k//2v3PpA9/zvW9gqN3OZ3SsnfHD2g/smCS98Xya2+DQaCMJOzVoLGsIaNKYt9FYhpIGW0U5mHcSrg2Z9J182Fvu1PcLGk1rhJ/2vRn25rYy+ODS6JiIXYa4doqwkk0fHAdG8MQZUpWR2f7FcxlpnCYW2Yw+MR2eLf1oKCfyZHc/S/n2dRCAZ3+3TgAVtngrR5gqV+uYY8mHlf0Ydzow9H0dR29GybTOzTuJR/6tcwP/5nFJYxybUV/dN/1GXYrC1PIKU/yV4em4Vb8RsMDz67jAHO0YeSDqfsL3eC/xQUNnFB7Y69e3oxv7rnuiJxFI1y9fG9h8OroWubiCU8fOJEmzcXtvhKKbelsXx8R4r0at68MERLHBXk6/+Ru/Pnzms58e/rcf+1+jb01YfQbK3/NM2Kajo6rLkS+lr/ODEYwpHZ+UXJcM5egSX6XKU2SAddZmEDMQ9q95mb4xcGmPY4U5EAdv4TvAKWEE4iqO02PrG3lUf+sznyOuZGvYw/FUy/1GihArBzZji4NXB5/OLZdyuTd7nHEa/pQHlkxn4ulNkyfnG4a9c9Q+8pL3Q6G+4bf1t8jtoqMOR9mzL77ERvj3x3mWsfJ9krmmPDXXrZdMpaUexNf66/mE+yQRV9brIDu2spYN8l2ydpWowM//8y8MX/jCl4YL528d7rnnHpZLupS3osXE34c7vPuB9wzf9e4HhusspTS67Dc/9VvDm2++OZw/fz6RZefO3ZoTK3VuZPyhJ5c6dC3v7OxEjh7ddo4pi5fj2ck2HVOV6j2q4z4OHPRaOa2Z81X2faXMOqSMMtI5Jt41nnfp6/hLZCTdWk/W90Vl7ps/6zt53/rse8vij165n7bbT7jIBj/OiUWZPt57mXq8+r5xpnFsF7Z5znuQ95zl4Bn8g0ZxXTBFq+saX5cbr/UmHVa+P6tvvaNuhrHcPDee5qnxOyaOvalhvG89eT/F4b1JWB5RH52kaX3jMfcPDeZN1+cr7xzmAHWJ7m6ZoIlT7PiFjY0TF+izXpgL/eR+vp018A1rYHaQfcOqmgFnDcwamDUwa2DWwKyBt48G6m/bKzjI9q5e2X35xZdeO/jug9dxSpzj43/tiMgAP9D7I1xjwLJJg+yIEwdd3uZf5OvbX9MUAwDjSWcA5hLGAs4eDH1xLPAkQiqg+ZnS8H5hENDqPSbHCLw0MKxoXsbGG7Juq/6Fx7qub2DLo90iwrQnUkWAkax+io4MsUpD1qVniXzDKFVcN9xfIRJEGTV2jeaSttc6G6RrNLk0Szy4ZkJnj33IXMang8x22zS6jhgPEwcnYGwTWYDK5WEd50YcZsDquDGiT/zH13GGECkkrGMRMxBADWjr3K/M0ch/I09ISnvrtQyx9KMdpOHH2+grcDXu8kV16LYu2wi3xTplKb1r1AaYutqHTf3E2Kd6OZ9qfuio0YG4p2OBjcfHALjg28FxdnCKyB707X5R5bQrPuLAQh5M9uJr7FhjK08a9kaLoI/IxphjZB7oCIKPffZ1unTp6vA3/+bfGP7En/jh4QMf+ECW2hl6sT/uoQdYcOtwMQJL3F7KY+SPqZdqcSd0HEbl0PBpYGzQSzkO7AuvwOmIGv3L6aPehIFYpp9OHaNK5NPx0KbO/Cz/NTpCascHPhxfeXIJaPO2eWJreOm1Yfjy40+z3HGLBaZAMZmcE3Kl0a3mVqAjWU8CROElEzTEU/KQxYFDPxhRbjHkWR+XPFKMjuyvfmv+6VC2AVhxhT/HDycP13H27frCo4/hIPsDkU9H2xHPg7yYdAgcsx9IpGdSD9ETFUFJWaegz6X7yAXOOnTszN/e2UVHq8NTzz4z/OZvfmq4/Mal4cOcTnrHnRfijN3k1MnMy4ybuMR/bLjO82d+jFNl3/v+9w/fxVLKT33qU8Nv/cZvDK+//vrw0Hd/9/DAQ+9lCSU6Rxbl0zHpWOzz7jz0QhebmxuZ8w4T26pn3st/PSOCl0Ot54qRd3kfwH2fgKvcjln6MC+NQENU3gE4w3gX+yxJ2z9CeK889ODqMYSec07lLcag+At9oVUmyQgofsktJV4rY2kp76cFXAAyh+Q3ex3SCVUkyYf0rM9zUghDR1q+N6wv5+DYiZ6BpR2UwKrXTMmxHwCZULTRZWQlbRIVb8thdGnRsaVSyuiktINufGPCh6kioHUs+kzCG3WNTzn6VMyaJvVc1nOktkz17x9Sh8fe+yuvB2XnRnw6x5KDSLz2VX+eZtqYogNLo858NwopnB2sZ6/PFXTn32z4p+dwfWVjuHXt2PFbaGANK2NdjkS3UeCfKzq1ssBrKqnrfv6dNXCzBmYH2c0amcuzBmYNzBqYNTBrYNbA210Di+9jP9b5XN5hmdtFbl7CQrybfK2WmLEAqz6sV9zjyailfKQDgCmxMCCEGeFSv7+/m3IMgPGDvu79mtckKOOAm4URYP+Gsd5knU4Nc+lqOFT/au9f65q+dV3uvOtuLr9VH+uE6z7S1YbSAI2BKC0aww/3uzv7WRZ4+fJl9iBjXzBsGI2sY+xh5Olym+snagkW9/J/AoNc+TeJ7rG8ulV61KDXQaQFFSfb5kGiULaJODtGvYcAyJtX9AC8RpzGsnXS7HZ5977lsDxNtmloFcxSX8JYV2M8jtWIR8dMdDHCqANTcNXtDfSsl8+l46gM7BE0WdHvOTHkVEAVuMLG+DoZdeAog3oP7cm4QHlBO3h09oTXcgpkllG2zqucY8xhnCXKrhtAnBuM60/+nZ9kDC8Pf/Lf+jez3xRsDwc4PW0vnDqsSp/WKZepeELvY51lk2Opc8KknuSldAEvqbGlkvhNPVZdbrq2iW25NK3gdYxleaQA3GePNQATxUXZPb7WTw7DF7/4teHipWvD3slTOKLgRx5x/EhvQSt6pVF9HypPOWcP93G+HkcPOm2J5tKBpWeilnw5gWSO3JP2cBzGWd57TOloaOlDk77Q2QdPItRw7KwA++jTL2SPtNOgaT0l56cdMs2noprkvXQv5LKsnuIYQ6c64HaYN1dxrj7+xJPDr/zqrw3nb711+MhHPjKcYSm0z0sO18Ah63PniZAOq1GkDomRYNK3fIA+jqPPD3/f78t+Yz/+4z8+/JN/8k+Gu+6+c3jXu96FYxGHCc4px9j3pPgOeF59Z/gsm3Rc9hzosbZe2byyzJm85WoZu73nVv0BomQWn/uOScfnc02HGbqpS+yd1MwyiUu8U37s07Qa0nKNoXpZtgtrahzi8VrSrvERpmEb3p72E0X3t80Ueup8lMFpQ23KdKl+VpFaT4VrOZertWC9F9fNMEWnouCASBfrTObK4lPXvKdtInPjFH56L5zzqvVreyfhrFem/JEFWOF9HTl+y7Tkp+lX39LDuNwyQPSHaRbrrhw7fn1n9+z68eO3fP8f+6Obv/GJ/6f5CtyUxyWd+W7WwNfXwHRGfn2ouWXWwKyBWQOzBmYNzBqYNfD20YDWQFkE9YW+gyH3Ah/3L2Lg7WARntKww1DgE7z+Mq7RoPG3krIGBMZcPr+1YozWoMyFHVXOGqIlsucNVPL3bwwEcfhNv5YNvYu85XbuqF7LftDbx1RL2awrI0/8qb/JsGkjwNzUtAJLnXj7EkZjxSTXgUWY4LB6pJF278OPvGEsj/J476mHbqCdPZXQ19HRbpYJXrt2bXjjjTdCQ1tLuu6z5bLLkydPQo9TGsm3tk7FEWR9os4gtbG5FcN8E7qOgZFkexiN13eINqOcfYhkzFAEZDC67ATON3lPdNG4J1D2AoJXpMq4eGfwBSMQed3bKPKO41t6FmXppfWn2h1X+8cRYO48kAdSVt/mrvWZgg2R234m8asH8QYj97AcHmy3Pvs1kTsfvORP/RIfk6WBOiycO8WNvSRT46djRKet1OyXiC1oyId1bl5v/8hvBA57Um1unRgeefjh4Wd/5qeHv/RX/vJwz733BkYdu4ecPBznlFDTHk4i9WuUjg5T5370B6x5UgSiPmThJ9U6LusZqg230Z/A6MPnIw47uFInjlVFtIAT2o6FLYW/8dkZeZQKAsHtM2wdDpJEv+DI2jx5Ytg4NQy//vBnhm2gD3CK0YFow9KfYxEGw0zR8PaI0MQVliUe7VIiku/ogH44srJWk7mFEiRViXuXcrq5vs61JHniPoa8D6vzadInm7TrBFZv7Nt18c3Lw2999qXhYx++A/7BLS304n/OOyN75JW3CffwP/Ib1Iy56B1XZ591LiHdJirw6vWd4dLlK8NnP/e54Utf+tLw4Q9+aHjowffGQa1efXZf53RK0+kz9RymwM/0GRCp+HV6OR/e+76Hho9//OPDX/+x/334ib/1N4fbzp0d/uAf/oE4ORxP4bxyiiXwRoTK9wq6DP+OMdFghv6Iz6R8h7wvlVk9Z2zSUrIFpqYQbb6n6p2Z6DHwORd83uvZqo6FY3wme6xHHUJkAVuOb5GP48eMU45K0JKl9I+GoV3jb8lnylK9K8ThWNUfUXz+lFc4MbMmMPk+uMQnXlO9W+reX6Nza1mzczIaGZ9lIO3HHHd8vO9LOonKJIeb0G1pGnOiTplfdIMPaDAHW5fCrBz5XNsuLuddzQNzL/sFLojHOmehiQAAIABJREFUAhU9V+LgpJyosvRxnAKcPCORZ8Q5q/zj+Du/2FfOaEGnQ8ki/eIj/I731uWkUyqzjx1HRfMeckbws3qCZeqnf/pn/sHWX/yv/8LwY3/tr8o0jDoeYX3+mTXwDWtgdpB9w6qaAWcNzBqYNTBrYNbArIG3iQb8wh+/8jHCjx279tBDDz3Nx/1T1F/lo/+28eOeT2u/6ssgUfa4rvxgx3jpE9WsN1UUy06MhnybUzfiSbtGRJwE9Jd8OUGKDeE0Nhre/lODLwje4qeMmTImps1N37qG6XZpdPuUnu1v1WZ943DJm3yu4oQ4JEqkIu3KEDrBfkbsA5PNvt2rSEPZE/Dcj+jKlSvDxYsXR93oqFiL02yDvba8jGZpB5qRZ+67pfw6FDSjdazpINPY0WDf390Jr5hI5VybyFS8jrqHNaOnHLkbZEbtLZP5tE26OloiZ4xKx3/UzcJ4rv7iNU37T/Ha1uOobuOkGnHqbGra5levXlW4wHsyYNNXjzo0DrbYU0tzEJLCF17lKidZ9jKb6EHaJumKS6NSD2f4Y/5ppP9fP/G3hh/4gR8Y/uBH/lBg1a+07OMlMfuapGdf6/rpEcY6DfBpagdA4G3A09iw5uVAQP7os5yVfXKq7dK07xLr0mi23WR78SSvuCrQDSyynxsORiLwXkedv/Olrwz7x5k7GSf4j0vD3jg0Rp7dvyoO1zgXpKncyKuzahVHwjFgcTzlVSBDMfTJ3WxfOJ2W4hIPKVzLoxcMtdxp5Cf7zOOw0+l4dLQ2/NQ/+KXhX/3efw94ngkiog72t4cj6GV80UPmAY671uU0l6yjI4zLHS9vXxuucYrsxVdfG77y2GPDs88+m/F95z33xYnl8/omTrlLb76R5/S2W86FP3XvPKs5Vc9Y+EWnRvhI07lr7ub8zpl//PM/N/zfP/ETOeny3exX1nxtbZ5IH51Px1bWg7fHFPLQw7GE4hIFqACT5Fw2tc5uzn1n6hSVT9+lLs2zzj3HTMX/6JzSEcMY1FV0bJdP63pe26/p2NZyWL8sL/kUtiN76bjAV/Clu+nzIHxHQApjObNEWs62lItWt7da+jmwXt57jOzTcnjfjjvhpqn5b7nFG1ckN+LOO8EOjFXhkTdw0+YLovCS+0CQproRp3OieQnA+KMjtzfSTzvzOdIqM1fzY5v3Jut7TKzvZL1lL9vNrWPceUwOD3WM63CGxDmCyc796z/8w8OP/dW/Bl4W1uKNK/jGNuezBn5vDcwOst9bRzPErIFZA7MGZg3MGpg18PbSgNaOF1/a3BzsX3/26Weevuuee5/GaL1mvEY5xVb5vj7k+90PeCIUgM29xr6dqWYXlPrgN0qFpUh+uPcFSD7m7XMc50Q7xzSqNerM12iDhqZ5rmwaPhoE1sdwKR9dGQbgFL98t9EgHZP1bTwUzyPs2CZMt3sf+JKE+pItuGmzv/fylToMeo1XlzF54p6RDHt71xMxYHtgY0zr1FrBwVV7Vd16221pWzh5MKiuc6LltWvbMfaMlnE51muvXRpeffX1wMqj/Y0q2zhxkn3Gyom2hiONTWWiu45kchwcGPUJMzWojEs78hRPfNGxQpLKSZWhB96xRZm5+BXGK44q+tGicei4WHBuTHVolIepDdTl8qFy8AR2YtRFr8BrgDK1dL3Ca43bAQ5AwlJwLqzHebGDPq9euR4H484eDjIdFJzW5+b7HVmkXM2P81EnUZJzgZvi3/GMmiKl+0PJ9s//ws8NL7/yyvAX/4f/Lk5Ko9W2if5zibDRZaU3nZKM+9pyX7nMSyNlwBZq6kt65J5OmM3uZcIHJuoRCl0C03COe/ilT80veAq/4kINZNNnwf4mR8TxyMykrxE5OmKcp7Y6D1aZL8P66vAbn3l8ePUKe7qdOQ+5olOsQqCfKZ5b53U5BMQhX8x9I85Q0qHzijEZ1umzR7sPrSn91e4IOzpo0oZsq8ccf3BTUbgdHKYVuswcUE841tg+afjcl58YfvofPTL8yB/50MBOcyNrPlOe4jkubw4m+o/j6zx07zH+B25luM7y5ivXidxkU/3X2Wfssa99LXv8fexjHx1O8Qx5CMFlTq+8+NIr8eOd5/TJU+xrJy86nvP86rTDuRYSyL5H/fWr14fTp08P6y5Z5dpn6a0O7T/wh/7g8PnPf2548amnh5/76b83/Mf/2X/Oc7o+nKCNpW6LOSleHWw+/86PCATTK3rK1P24d2HJwXPsRCUxkvz2s2aUapmsaBs87DlIq7wHpWPhMPmOpd1pFgcNjZmTeb4Kb8Z3HMLwI7Ebks8Tw8w4VZIGWJmsDZ8xlQgpm2B5g9Lsw95Y5PDIu0h4YzbF56mSxW/xVCe+KoscV8rzxHNlsk+Pi/i8nKeBH+d8nhtgpauT17wdhY1TUauPcNJzvjB7RsdW9vmLHukBj8J6Cauu6l1ZMlBBffXPY2AhlfAHXvt1iqyipM53quUD5oBPr5gdMiSixByGn9o7sHGUvPYRylSPXenQsnx5GZmcaDixHa2e2b6+eyvL/jcB2UZOFTaOVI9/j6tY5jRr4K01MDvI3lovc+2sgVkDswZmDcwamDXw9tVAfXXHrDrQHNh717vufwGL8xk2fn7DzaRN5fzgg55PbDftrx2B+diPs8iPe1MbcRrEfqQ36v7Yr3xpPPQHei05EkOMkhHbv9BfA0OcI94ldntWsr2Mia4pI8ZSGTtlWAnThl9ojri7fxla5Rizzku4zuPUwwDUwtYoN9JInGswtbpR0QRGfwWPUTw4FzR07W8ydymghp8Gsyfk7WPYa+i4f5mRZva1zftsFH7lGqvOcM6AS0PbSAwNdE/eO3GCfcwwfk9s3hb8mFFFC3IucWvep/RbbtAEttusl7YGuktpp0kZ9/fEpyzTluUYN55p65S+OJq2sJZN5tI15eQ/DGRPOFxf31xEcqkP054HGqzhrMoywKUxGzq0m4/2ZN3bCVqp14BEPyb1/+orF4ef/9l/MPypj/+p4V6WViIdfGgAs08Z9OVLPjXaM47gRoI4eCIrpOKEdNnhmCIHlqz07FfKqqdEEOu9XBelU2uRGMNOjq/Re0CnKjzAUzsiHZ/Q7w5CBid9wKmfyqVvR1g4n/ztR/BAn8xpkYSBFT5xiUP+APa5Di3mtE4O70FHMBeGd+Y6iHBKRhZAbYvDS/6JIMvpl/KrapFD3pyrraMQrU65JVq1xpv+WWYGjqPjm8NP/fyvDh/+nvcP7ziHgxTHqY6ORKbBrwdVHBBt1ik6YX6rRx0Zuzg0XU55Fefmi6++Ojz9zLNZ+vmhD31ouPWs+5YfDE9R99hjTwzvuOfe4c7bLxCtqQ+hHA3BBx3nWfaqA7fPj/1Mbsp/G47uxZzl2T5z9tzw0Ps/MLzywvPDwyzT/epXvzp8iM3/1WfGH3wV6bV0lokvDsxxzmc+oPY8d6Ne5CVzb/FevfEdFIb4sS9o6p2ArioSynlS9JxS5bS2rt5hxb/OF+vaYVK4pOvVsOEt/cb3LzSbt+bBXDhT92+dWZu2kXY5nCbPe3gYcUPX6ZPpN/IhTqCjw7qv3ym9vu+8x6fKKIAkX5263jo0kOrua973Lafv+JsjPxtO56yYhaXnoq+OLGEaR9PuvHRf74csgw+W0ot9wJj+zUvncWKHVr0v828ROvS5UG6XhzJ/Tx07deLOu++++wJcPAumfd4bhpFJXoGXyrBmTrMGvo4Glm+HrwMwV88amDUwa2DWwKyBWQOzBt6eGtCaZ7XP3s7wO5/+9P/L3psFe5Jc93nVd++9e6Z79h0DDGYIgCBWriIJUoRkiSEpFLIjFLbCEYrQs+wn68EOy69+kZeQGKZN0SFaIVsiJVG0SJmgRBIkQIIEAYJYZh/M1j299/R67+27+Pt+p87//rtnAOqZU9ldt6oyT548efJU3Tq/ezLTj/oLfGS/nY9+PvL7Y94P8C2dxvHj33yvc3jtodPhBzz1KvlRvuecJXomUQQ6EIAOHMbgmKyTxbX5frdtDwGGOExGW9C2yXwa0Q9PnZbT+i2reXEYyDPfox0naSwPn3AsPqGBp3BW89SBMmqi75vXWC35bCIWx9S/4u8naufwgcMpFsiyTZ2Yw0Sp7GcnvOWVxRxe72eq4LHjR4aT954Y7mGh75P33jPcddex4dixI8P+gyzsT7nrk7mgv4Cbzq9tJAFk3GD3S3fAvAAY4FpnG4yfNC2rAOZ8Mj++nuhJdP5OPRiKEz1Hv3tOmrpW56XDiv5RF6Z5vfa1bZmkqWvbLD2ar7MmCCGwIuBmim5pI871yFsQ0Cmn2oWA0S3WYoudUd8opE7uVtfOt/VrvS/6R5SjxxJjoGypS9SOelOuX/mVXxmefOoDw9/5O38nEULqz4X63XXU6D1lss5iAIcCdeCYiCXXiTLqL2tJYSdbyG6ZAJVRKK0D+32nvhPJBZk0youWaAM6HiYdcvOt1TwanJNGgE6ZTFVeUZ2946xl9nVplbW93h6GF147C/iEDncAoeRqdA5ijg6zTAKW0dmSPZz5QT9sZZGF6wtxox7jFWDYaLIAtq5L5jhi59omvDrJvyKgChRNvm2o0/FZtl/KpD52lvcPr565Mvzj/+eXh8vrbE4Bq44Uc9p2gAqY1PiWfrMTKfozsvAaUV6XLl8Z3jp3fnj9tTcydh/98IcBx45FT6dPnxm+9rWvD8ePH2edufvzXNFsxsyx83C6p/3utee0qfxBgP4aWegagJuMedu59vno44+xftkRohzfHr7whS+mrX5Os4slc0ndwVWbdGwytqjS91/zIbOeB/on+NnP1t7zo/aoND635meMAYlXV5h+jcyC5NoGIxE62zNa1zp7/LijHx3hpTwtk2cGEFFKRm6Sutz2lOCd0yQddhRJqbQd8ZV+8g4UKK2+7vFzDHscK1ce4/sGkX2OZNnPgmUepu5LXSuR7/c6m3d7Uq46rC6cVb/D6hmKfnnmZlToNfzVG4fXHj1O/q6TR8tTb66iiwpoLf3AbmQR/sruO47nrv64YGtF5zu1bhw5pkiqe8ay63k2dd95i0ElH8Tz+UTf/J4BF1twEnTqASiv3by5/sCN9Y37eV7X1I1sYUOt/LYOz+nHpIE/TQM+VVOaNDBpYNLApIFJA5MGJg28NzWwSwQZzszv/e7vDFfevvw208vO4tTcHD/MF/kQX5h3fPww7ySNDoTObpz9Oz7q4zDEySiHof5iXo6WDkA7A81HvmO7acK22lEww2vb63rmNX3nNX3L2eVd37Op8/tsni6EaT6vcvYcnvl2NnGqpV1watPYdx1np0Y2SNZ66Xv5LeN0L7JTo860xxKOruuXHTh0MICY65E1H3fX81odF/1S7s3z3nx5t66Uw/WUTK0D8wS6lDXXo6ytS2nN914X1et5Z7j1cee5+VvPsi63vteem7fX0pvvWb0ImvZ9zMoBIAJHO7FfpkUdTJzJONVENMmnnP+9cWoeKRvbNs+jk212+1/83S8Mzz//7PC3/tZ/zlTOg6xJdWX4d7/6a8OXvvSlrAU3axsZ5vtg/e6H5+bfNHe2WfosCaS5877bsV540M8ZwDfKb79NLXvaHQ3VvHmejp68ltYWh1dOXR1OX77OFMlVHPvbk6AWhA56wAhLlcVpwzryOuyJ3qJ8H2BYplhaJhDmkOKgx/En0k4QKTYuT65Nrl2mbJUqj4zq49jX1LF9+CrK4oEjw29/+U+G3/mjbwyb+5BZ554C+cip9ZexB/gM2EHZDRfjv3KNaZVXhlOn38rU2A996EOzcXz77atMhfz6cP/99w4PPghuMNqqfJXBKFCPtENeg2SqODpBRiMKL1++HF0JoPk+NO8udsW85557AFXXhhefZ6038uXZfc9YjX2w3eanXtpWOm9mA2OZwJrgUtEBeCFHvz/BxuDlaHveeydKY6p2bx91+XRqutaF+d+pfJ626Yr/3vNtn/t3hDSWq4PmWX0Yx1IdjzSeLes25uln4yERqWn6XLl7cs/nd3tNM38OXxAtaex//nCDvF3fs0fL0vl38phT57vSRwafEwgF0Lo/nuXZuu/25D/fZuqNMlrWdZres9nQ+eCVDPuGNUC2B27d2n5wxcUw95LGUsaxlzddTRr4jhrgzyBTmjQwaWDSwKSBSQOTBiYNvMc0gJOZiBL+3m0Eyr/+pX8xPPvCizd/9uf+8Rm+4c/yAf8w5yUWtfaP1MYmuM/XOz6y8/HPH6l19NrRVJOLocap05mzPocf/UuJGipnTVdJIMb8/vC37vjx7yVlNulRDl/TejbN1+t7y5TZMh0SU9M3jdFScqVzKdvhz/7hbTQE/Vmw3O6O8qXMazrkToobm+4wuZF2pBEo0GkVtDIZdWIdI6DUjetreS8wZkqEBICP8QOmOEw4VEvj1MIFFitfhh43PvWNLggd3SYbepaFAohbYXc8ATcd+orOah1LZ1TYqF8rkDraaryNTCngh/JVUmelP2Eqdym0H2AZMoBQh90bU+t5bwpcspUd2kzng63RDOoz/RzbiX5wrtWP+fbH5OYH5qV/5Em3se6GB+vD0cP7sZmaAmlEjEBJjVOqhlaHfYFpcKYGGap0GM6cPj38+uf+3fDRj35kOHj40PC//sOfGX71//214aWXXhoef/xxptKdHB7jvMI4ynd+4X9ldMpVpl1hA8rlIvvm26b6xpIpr9aSR5l8jHiyQBr7pgoS4YH88pFHyYp6oSyaeq4ENx3f8EHfop2JArPvyMG0aAAKF6nfBmQFXGX24FeffWG4vo1tA94sLAJk+fikUU6OoX0JL64TfYgcaQO9cZE1pKTBtraNUVlG9n1MdZVIPkaU+XCPcsEsSRk7FdjHXeiRZbQHy8t+KrpKHrtMtVxaPTr80m/87nDfvXcP3/fwcfYuRQ707XS2RB06HvDwULdGFr599fpw+q1zw6VrV4hYWhqefvrp4eTJEyk/f/7C8OWvfCV0jz78cDa6UK8lY+04qWLRpkJGf5abshsh54Vl5CYSzHUDBVIPHzyS9oeFrdinQLVg1nmm7J4/f2545JFHeA8ynqhHGdWXYOMC9JUY50Ty1Zg79oI0/X70PuOMTvL80OdF+qUNCIzJS1BMORd5R8QwkF1abpQ4Z4dufizK1qqf2lradTzg73UGkp/9vi17tGxvPCme8ex629vs5Jt3W9E5/KXDsusZP2T0XaCNq+s92RxP35OONeOLTZsUSbk8Sl7zlSfFdDVPWsyx6Ass7nJHVYnq557czhp2owan526xxl1+sdG2QLw21rqJTY7tp69pmyg0GdAH++i4GS1m8sk3LY/vOQ0AbvXOhP8WwuR3Au26OUO/P32nGk1N7xXWLqInLqjTYyDfhjvz+qENNph2zEOaacHog8dklWno9508efI+fhe7o4kdlyk/fK5toPQrzylNGvhOGvAtMqVJA5MGJg1MGpg0MGlg0sB7UQP5Yi7HYN/w3De/dvP06TdP8fF/CmXcVCFO4+C0Sx6+iuR+buvM8FHPgcuTPH90eWfsOUHWEbjxw94a5aR2eRyQkXfXbX7Ns2m73PzO6+u+v7PufJ2+vpOmeXR7nvvoOs0/UQdkdh2dpSyUPjqe0pfDWrqav9c5u0nUi1P9jEbJmQgW1z9qh9h25ClA5NkIsT7MWwYUM7nxgXCeNGg0eag5qcGJlsNM+Xaf+uxoeFjW/etzcaqf0nSd5tM8+77rSVc6odbYF/NMytPHXl7lN7hoZJ71tZP97OaZtaHQbUARQAfrOx3MpD2ZWrZu27yZs+sNCRcy4Jj6W1lbHf7+3//7w8/93M8P11ncnV1cMxa//K9/ZXjllVezK1zLV7VH+3a6FHJ1e5bNR8+Y33qwrHmYp9yOY+f1ucpGAAUP2BZM5kvj0dcpGH+YZ2o+6s/F3Dfwpr/w5T8G1DqEn017cAxLyJ325jpgMCwuI/Bqq60v+caBp6+RBoAt0WWiPvHo4Wc9WYzyIWXAupk85NPhHK6JJkBjhdv7U3aOUpCTNZTQ65krN4dvvfrmuOtm9S3vDGSqsdaOBCp2Ez12kciuG0wxxiKGBx56KOCYtmPSXpym69iurqKbMpVZmePWu8teIQpN0GTbaZHoz7bkI41ngTB3WfXed5n9cLdKMcItnt+DRw6jW4AnoAxRC8fa5Fk5ug+dZ36XhZAfPc6l/+qv9ZxCuTxGijU41mPffOf7Ns9v/to60pvaZvpsXrfbvC2bP6QxzefZt763P9btc/Oxzvy1952s2+CSY+h9dOOZo1Pne/9uvMyTxhRarnsqtn9cqDxlY0woE6wSXPcPHUYhsrA99GWyYXLHjzwt1LMdn39lNHW73Xbnz1fvsj47BgKHd45F15nvn3XmD2n6Xjp4RLSxzhp87zl44NA9RHEWQFYV6uGDfkqTBv5jNDBFkP3HaGmimTQwaWDSwKSBSQOTBv5saWD0JegUQTA4ffZud2l9a3P7DbzNN4js+gCu3UHdAL6rOc15l9LqIPQH9/jX/GUcXaZ35AM+ZflL+AiGQYNfQZ1yLHIDj+yamDbKiZl3OHQgdEeMvjHootPoGORWmnbI2gGxvPl0nT53mQ52O9LJQyz84yRBJvnKzzIT7ho/qy/2zagOwao4iJQtEQHT6TYnSdlxxBLlRX83iI6y3LWTbM/olNwTjabzvRkHXMdHB//WLCItbaNPF4ZfZNqcu8DtyEOpwDDLcaferO/wRn4ZOdQ68srRfaa3VR4Oo2Noo8hkj43O8rytjPIhORrELGRoFxlHgQTL1IG0Hk43zb1T9dQdR+mxQAvbNV+O9nubgcVsQhMgBUDMaDX7I0fXYGtQSb7a186q0SK2Zvdsr0CIjOPY/4BM2hxJXjuAkb/HOlEvEin26GMPD88998LwNqDIPffeO5xgAfZLly6wllatHfcVoo6OHTs2nDhxguiOcvgFhBLJFLtA/oyr/MuBda84I2ECkrS+oI3ZlhjIWraqTG1Xqt9rI0SECjR0OKoQyUpXdFW4cGSTvDwbkQ3SKB6bdDrk0urw6qmN4eJVQCMW6DcCDEuXUVoQLAtrh9o8Ktuu1zu0Lf4V+5WI4h0X9/eBgA+KFpUlkwIJTQJf8uG8FyGmVcpbiYn0InxmEXCNkY/9ag/ZAKDrLvD8YKCuSuauh9c3mPZIRJzP3DLtabdbRLmWTRRb7eDs+cusHQbwzhTlQ0R6PfnEo3lems5+vO/xxxM5htCxffVmNNjpM2eGbzL18rVvvz6cZy0/o0E//qlPDj/64z8WMGwJuo3Nm9jfakC0BWxjm400NjfXU142ujlcJYINpGV46oPPDIeOHgmYW9GCytkjVtfeC1wLYmqa2ox/NEBTSRlT882xjOfavHp+fOe4G/D4jPIukH1shtrqSDpg5BrXkacNpd2w3HufOd4lz16eVdxt0n8L4ws3tmU+fPMStlFa8f0QO+E6dgRF84wtofvOD1/7lTa7t/JBdZoK/S22JZORgVVqv0p+aUy+A0zyysG1NJ3UZgNiAmBWmwfalJn/1HGTlVvYT/2+0p5Wl7eHI6wZmWmr1HMcZOE7Vfvx15njIQ9/b6V/Y9M+n/7LGErPEbmyOQa6kY6xCK8eE/MoN/qYqpU4K592Uf2qBmxb0Nrf1faxNmGBG4moQl+IMluhzokzZ87cvbO1xS8kQW/lANLdwUjpw5QmDfzHaEBrmtKkgUkDkwYmDUwamDQwaeA9qAHdtLi7fES7U+D29cOHD768vLz6Mh/61+ecMz6vcTNGR0QHQeegN5Bv0EXnpafwCRR0aqfBOqb5c/iM+dKV07VHI32313VbDu9N8pjP815ZOq/bK+pyqLpv5jWdTkinOEH0t+t67gW3vbaO5/m+ee9hUifzbSjPBgvNm3T9pdOR3yBy7CbOea+F5NmIKZ14z9J4NhnhYrvzbbsu0dI+o2MEGPbKUyHOUemhdWi73V9plLb5pc7cffflzjrtlIuR6PBb3rTdjrxaN143TdN51llsHVnPtdfcnOAWUR1G8vSaS0bvbKEDQQynvpUO5Lonu3w8TPLuPvY4njtzdvijP/rD4b777xneeOMNFly/NfzgD/7g8NnPfnZ4+plnAMruH44Cih06dATb2R1eIors5iagJUCAIEFPH9aRdkzk65i2nbUOu13l6Ovue8s2f/YaTgitj4v8nFtHlt2Z5Bm+jK125GGy7j5AnF3WxnoB0OfK+iZgHdNTcZJnKfwZK8/Nh0Id7/A0TyfcCkYpCnIKiBk5xrWL8wfNFAw232c85WXzMJo15YVRY7SW/rSe5sdGelQdUGvWL+oJiq6s1FRCWQaYgM5nyvou7H8LZOU6z4gL7Fv3vvvuC3AlgGByOu6NG+vhbR3B7NgRY+fGFp/73OeGZ59/frh242o2aTjCYvuf//znhz/40pfTRtdxrLuekY2+1wJuYxfahFFla0SPPfXUU7w+yzZt3/oegrum6DdX4/sMPtpV53f/y47FI0uXzUOgo3neruVqS9az8rFteZoX2+DcbY1i5NR1Ok9dtyyWzZLAbWxmL6+fLWmaT2x4vO98z52ad993G/O6sEzeAlxN732nbst7yzt1PwNGkSldyyggljZ4HniiA4wJxG2wKcSN65tsfHIr9nSD58bn3+Z8tuTfPGyn2265+37W9qjnzreOZfM85GkU4jyP7ofn+TbrXi72Vfh4zy6o7xpkKcJOaYI/vGxsHDty7Phd3/8jf26/z6zgIDRW2hs4a0xp0sB30cDcb43vQjUVTRqYNDBpYNLApIFJA5MG/uxpwK9rP6H9HsID2r556vQb32Y60is4dtd1nLNeDhtd8nFOsNO4KD0f/Fmk23VW+ND3w5yLuOrtGMzW8MGPHj/ic47LPOeEWZb6CNDneXqvddLn86Trdt6tTuc5XPP8+755eW9qfl4LMhkBgm+fY562nSBBDB1nARsx2H+ZAAAgAElEQVRVF+erHJHw0pF3ulucY3QoSOEhMNFAi3WWnLqmE4P6bMcyo1ausiue0/48rl27QVs7AcyU06NlSjtEDGVqnaAHY2FZl+MdBYRyjBxewYgCtMo5sz+OW/WLPBzSctwYE/XCQTHJ+l5DK17i+NOOyT42H5EMyQW+BDFqp8ragXNp1c0FlgNUWMfdJXsM0z5tnyRiyx098V6jW3fxNFJPgELdbI7rvlmvdeHZpF2VbQHfAX7pEurgWr4NsOGi/AJ7Z86eBXxYGv7iX/ip4Qd+8NNZM0qH+eLbl4d1ovuu3bieXRlffvnl4eyZ84keunGjxmBDcGw8jDzBJR35F1DWslQkItL4/CBr6aoesQjLj9afOmvAUaDM8dG+SvtcChIgf8ZOo6SXTkdUZg8pLTMqaYmdVHfAY1587XX0j90xWPtYMN9plQxSD2YivRBMIWbXGasR7JJX1i1zsB0nIrQGQTGBMmxWI5B+ATAuYJu8OOwrhYm6CW9BagNXAI6UPBs/oLNcK5MgAf3bIpJHfWgHR48cGh68796sy2Q04jJtuT6XkVMr1NEepLsJ2HydqXHXAKiWeQaOHz8GDbpG+RtEoL387deGSxffDqhm9GaeRWTwuf3iF78IwLYxPPn+J4ZPYwMf/sjTwwMP3jc8wI6yf/jlLyWacHuH6CLsaJF+3wBs81nvZzdTn5HB59IdND/28U8OH3j/+4IXCjCZShe+W2pKpvcesXWvGbnZ7pPw4j/lVq53WwPsaDrvJOsJmkkjrc92yG2MFP4+f2M7sUV05jMgyNs0ntW1dCb5mvZ4CbTTKuXSzR+OrUmwU6C4cJeyc/lU3+Q9KgFa65u6PSOvPHxGtN8utz/dln94qfyi6/UX5/nAmdu8VZGqdNvPX7clvfbgKyKy8q6WZusWB2ef4Q0iSz2c6q5tOOau5RfuvESUQyDNNdKMdsszD18jvBL9R1/SHrrWALyOLhxHn2VlsD/2Vzl8tgE7Oz+A+EhnXYs9qv9S3TEOVhUcH/VlW0QaV8/oE5tHrB46eOToz/7czx38K//Z39AAm9neoMh2SpMGvosG6kn/LgRT0aSBSQOTBiYNTBqYNDBp4M+oBvho5gOaZdg58H4BKU6ePL+0vHiKj/Wr9lmHgo/1+Av5gNe5qbyZSsw3z7MpDoFOwXi08+TZ1HTNr+tL33khfJcflsunZfDeZN2W4d14NF2zbBrP8rN+8/nTzhU5xNo1ACdvX71GtFNFE8liBhjBpJ1c+ZtvW4JZvUujedJ0e8qvg5Z1ydY3ct1OG50bQSIjHGq9svn+6mzf2QfbS96o13YkzbeuR+tNGc3v1PfmzV93HUm7Pe1GutkBr+rXTqa3La8sDq++8tLw5qnXE61z+PDhbiZn+djPI8cODw+xjpRzNy+eP88aT2sEMrkOWW/IpmNrlGLZkPU85uVumebLjBh668yp4SzgmNFJH/3oRzOd0kXXv/ncs8Nv/dbnAdBeHO46fiJg0ltvnQkI4M6FRv0pm0+JPFtvyRv1N2t/jPJpGexcX1vPVKBZjbl6s1z9BlwcdR3C0NZ4yL/5tMMcTDu4dtFEPoCgW9y+8uZbBWg5SMgUy/baw6Qzz3XWI8MGdd5DJyAA3CAA5xRkjHZGmxXix8ixfQBx0ghyBLwYwQH5RE6cdy7SVH54z+FGFT47lceZaZOhAznYNmoQgPJxgKpH7r8bEWsKtPzsf54lzrvw8N5pta7lJ4C8emB/RXlhG47LpStvJ3rMdcGs5zNnHfVs9ODrb745vO/JJ4fDRI0tE1l2F4v6P8r0THekXGIlfO2lx8vn0WufVe3Wa8H/HWS/evntYYUpwZ/+9KfTvrJ6hIaz7dl+ZHeMSS2HZV2uvc/yMQ1xyb73jJIAIotvmPDDup0EpLptsSnlq3pFJ23rsc/Wlcb7Tr4f3i1VnfojhX3rMRxN+jYe8uy25dXXnd/33c78fWQf5Un04SifbUrX5647rwPzlNODESqS8Y8XaAHzM88/EtBneAUcG5/t4gMNFE6dDQ/aTPTVnErMNynL/LX3AqPzfZmnU25BOc/Wa7quF6b8sNzUvHMz+2G9umke0o91mN2MtKN8nA8vLi4f/tEf/XEq5FkfFTJjNl1MGviuGuDNP6VJA5MGJg1MGpg0MGlg0sB7VQP5KMer0TtaGF5++cXhmY983xU+uK/rMugw8sm+j7+WEyxCDh/lnrPLHVXGb/p89FvmR7pHOy8zJwDuxryM3l8iV6Tpj/p5+ttGgk97nQ+dcXlJ79ljPvV987Osr7ueeX3dZZ0HcejtQ9FU/QWigDrFMTSKhmQUycGDB4fn/ujrw5XrN4a7jx0djhDFctddJ9hFcC2gjvT8RX/U2e7Mid7ZWc1aZDrzTiVbWDjADnlE59k/HG/rCSYsbKH7FZwv9BwnW73yz7J9OOxQR52WtdxZT04+6gdQYqYXnXropTV1lEfr0/qmigqxTatTP3l7fAT3rJP2KNu3yODgVBrnAppCRumY2gQbLQ9/+JU/HP6X/+kfDGdOvRFA5EPf94nh7/7d/3q4/4EHEhHmtDX5rRK91Auq/86vf274lV/55eFDH/3eTLu8+/hd7BB4PlE8NzaI9IheC9DrvrdMCtBjrE1dJjLsN37jN4aXXnwl+YJtz77w/PDCyy8VmHKJaD2m4j3+2Psynpa7cLt8rO8UWC6G/SNAYVSTST2oA3dB9dxT4JTDSCmyyd+bfkp2+pnK/KhxkReE0V/pMfdjubwy+urUioyn/0oCxoBy+RrNZVzWNrZ65caQ9cf2uZWlgFYnBTLRVippDUFi5A1HwLWB3Sp91iKDoBeRLZp/2YFrmTF90Z0xBbwo2AM0yI8gJZkcHP8FeO4k0oi2wOCNNjM6SL2oW9fT29nahKf1saDl3eEHvu/p4eGTB4flW9fE7GKHgmFGkakzn7udzXpGjOhyKqVU2QQAHoLH6zc386y5jlyeG7qyCEgm8Pztb387dnSLPtx//73DdQDuu1iD7jKg2I3165FrmXXHnILrc+jY2o5j0YdymPf6668O3/M93zM8wxRdbT+L/FPH8rwfOasr+0r8Lfmj6lUPN2TnsO5iovKkLR06Dq7pqK7sg+/OshkrU90xUOc8fz66lrHfcGSsazIBOZ2URyn59Xw3jzy/CmSpZ2XzWrbJBggTTLINbYv6WffKW5LTEO2XfAQPR8OhZI6ndzCUrnIlg4GyUs882YXlyKtkr0aqbQikof1aT6veRd6nDyoxqfJjNLRhtNeunaHciFZMKJFhRoC5vp0RcGLAvreiG4Fk6skz487vvX1cZ3fRCFq/F3y2Ixd5ypomHJ/oieZ8bkjGoKWc6+abgrn7jCv1pHO8Pfe41HiV1qyvDk2253s8uqe4bbRkKRvlOWOx/p1D/LFrcXFtlUdinY5RE/6+Q6Y0aeBP00B9JfxpVFP5pIFJA5MGJg1MGpg0MGngz64GnMmzsG9pZWtt/6HhIx/+3pMLC4sfZ+e6D7KtvV/p+NJuYI8LjQPox7lAgR/lfHXHAahFtHUuGmDyI55phNQSZHN60Owjn3rW7RQ+o6PQ+ToKcQyk9Zt+JO9yz12v+fTZdqzbNJ3vuevPOx25HvsRZw86ncTQ0rbltp/2pMPZEqRxytna2sFMw7pw7sLw7ddeA2B8eTh37lyc8KyZRVWdS6f1qatlom/k5VQxk/kdSRY5KNuB9zrTxGxvQUHQI/hkIsp0LPF2UlftLwEsPcBC82tMYURQWVeyLrrv+1oPiiIybIfiJNtIP+s2/lPfF12Nr0PQqeuHDj4ZVwZJMNE8HT/Bseee+9bw3/93/y0gBsAD9iJEd/at08Nv/fbnhw984KnhwQcfyBpOcQrpi0ld/CZT4F566eXhh//cDw/HARzt8WWiddZZc2oF/e0/CADJtEt6kvaUJ0M0dkobFYwREPmTr30N+RaHxx57bHiV8XmL9l8niuj06dPDqVOnGEejJk9k6iSLWw+vvvpq6n3yk58C5DwAaLc/MqmY6udoB9Fh6c5Fve33/GFf+l75ongzO2lESdbDXgOAmFF8dnjsrD+qpUj5ObNtHWZYIFXoFtHLvtVDw+lrW8Ov/c6XhvXFg2BZbiIBEXwie7ggi3yRWbuKgXj2widcWbRXxlAJS3br4DJJl8yRVn5WFYTJQ8pl2JvJmGCr6r4ANWgyThAAAme8AOC00F1AIB+qk0cPDH/1M58c7ju4MKyyJuIyPMKJPthdxbatW9S/cPkqoNYNpiRvDwcPHxiOHT2UPl65dhMw9WIiBNdWV4b9gNXKZj8EtV5j+qnjb/6BAwcBZlewrUvD17/+zeGFF14cPvbJTwxPPPFEIhfVv3W0zwYuVoxGQ4qbTH/+8h/+wfDx7/0oUzMfGFYAJPMcoyPbEpSZH3+Bk9IlPaAzLri/CK3/1HV2qYzWxnI7bP+r0+mDumqezT8gEJSmgDec5dlArnemBt5yk3v5V+o2whv9MkJYowNt3ZJbcMzkmPJ/luxL6kOa67G96GCuDyUFHLs/aSUmEb24S6rJtgWtZjtQaijmqdPwKx2YZxt5dkaa8VSRjVRj1K05o3Pdug12q1znDwzrTJl1nUP/afY+w077XgWAXfLdjMCZEmxDJOWfH1e5K4/j2rbRfYseWy+pOWS3zEzZddx9P3JeEhSlXccybYw2U9fJmo13l9ultqX0ruokfIyRWIpdLCxeXFta+WN09vK/+Of/bH1z/QYNqCwOfhbn6eekge+sgQkg+866mUomDUwamDQwaWDSwKSBP/Ma0FHS+zXmaGH7uW98a/iDL3/l2H/6N//mhza3dx4jKoGt8Pzkd99CVh4jJADHIEuT+YFuhIOOSRxxHKdbOB/zDoNT5HTO9K3r433v+zwOBo7EnjNVyi5HqB0uJTNfZ6jqlmNU13FGykm4zZmQZv7outVC9cjrWf0usDMkQRmvEtkB/8olnwtJ8NEDqghcrbB4+dG73PXwZPhdu3p1+MY3vjF861vfYrH3V4a3zp0dLjPta9NoGvwTAQOdJB1qo0R0yg4QuXSYRerdDVPwzMgFI8Vujd6oAKTARfISdaOjys5rgAD3jwBZqakAytIO/aMnqi06LILcp5Pjj9ZndCShHWxdM6aJ9Bn1YhXpXAPHcVIvdV/t4L0FnHDHv/+ZyLGd7U3osA92KjSIQV6CC7/5m785HGEK3D333jdcIXpnnbwV1ii7++4T2WnytRdfos4+1oj6IayTSC6ivAQyjCBaZgH5A0T5uLaYbetb9zgpl3lbOL/Pfuu5gFwf/OBTw+NPPM5i3NeGL/zu71CP6CB2AHXXSh3+y5cuDufOvDVcIZpI0OTHf/wzw73o1IXbBSDTZ8cNHZQeAToBfbVr1RQZ7Bv35Gbsyt9XlgIi9E1Vv4fPQfOJrqPFaFJmacepmKY8M+TZhinDw9mWkhfvHntZXh0WD68Nv/etV4cvfv35YRewbGuwf/BVTg7BlCy6HyHgb10OwYkAWeRDmXunUBI2WnrNM1rt71OA1OdH+i8f2hA0sQseJs41nbQyUzsgi/zh7RMmeKdeUrg5fPxDTwx/6Yc/NBweNof9sF2EXkrXITMSyXpomTWjWGifXTovvn1lePva9URrGonpgvlnzl7AvjaI4lxlPbPDeb4cl6wXduMm64ltDG+++cZwERD74rnzwykAs5ewtddee4O1yD40/MRP/mSm4aK4RBjaB03/JmvTmQ5mE4et4XXA1rexxx/5oR/O1Mtlnluf5SVA84o6pZ/ocMFIJHUvE1KmV9MfARJ13mvx0a3YuX+p6Gg5x7eu67nxjw25hxVVSWVTyfOWVDbhWbuLlfATBau/0Y763O/Z+ee/pPS9HnbjsJrr+wb7TwH9kTthT/ZN9jNe4/PnM698vuNM2rHJKDsraDJhwtlx1UyhCi/NJNGR0PrOMwlW+Xulnrn0yGbpEz+o69vaseItlPGyju8a2aJFS2M3NwE8jQ40ytB3fDEBmM+mEAsAlfVODn4cu5uRpI+uIWafldnGw4N7+5f3oWNt26UASHiP+wePLP5PNGDeG4Jj2IV1lJkKgqVtIz0+nl2QLEOZHvg0FP/0mOLRrHbGCDRwPp7lfQtX0O+3Xnv12y//01/4J1d32Zrafo411diUJg18Vw3UU/tdSabCSQOTBiYNTBqYNDBpYNLAn2kN+E2Pj0FEBx/YLz77retX3r765urBI6cBEw7j1KzpCOAShA5HZd+S4AJf53uOQDkwftTryAgAmeY/+vu+6/R9n9tRm7/3r+x35lveIJzXcSS8IJUTpfMZDy33VVJ0LU/neTZPR2NWpmNC6r6Uo7JHp6uRKCW8ECPjVtdwipcPA6g4xfJYosdOnT4znBZ0uXJtMDLprdOuf/VSpmAKvpyAzjWNnFboWlBGRCUChWt2Eg044xpZFy5dinO1w9i4QHzi0PSGABd2t9GNIANJ2QOm0O/WTfen9INrRb9K7upfl1u/9eZ19Xf0o+5wp9Rr8/dMo6FvRxjF5/6FF14YXiIi5+D+FRZQv3t44OjhABmvvvTicPO6OwzeGH7mZ/7R8F+yDtCT73vfcIONCd5kGuZjjz4+/O2//beHL3/1j4cvfOELw0//tW8PDzz0YMC0NcCx9RvXhs2bq8PVq9fps1NYifpAd6urNd72yUiNc0T0GUF2L+tKKed1psH+6I//BONxZfj93//icPnqlYBNgpuO28MPPUrk0PuyG+GJEydiP65d1SlRe+hPwFfgqKfOWW70CWqg395B6U6KHQFmzjg2ln6nVGNUtAWO7TnM1p8vl4d9yhRJ1yHjmd2mbQNfvvrsc8MG5pGFvp0SqWfMkysuEdBEIT32BEYPtGWegATATdAL7UrnHVvz3wLryO24wBntLXDsADJahb07+CGaxY1TJTk7/a9tq8/KTGak8cxN7qkAv1tEcu0On/jw+4cjTCleo2/7Yt+CA4IcjrPTDZEJ/plmybXvJN8ztuF05Y2Nm8M6tnVz/SZA1iH6SBlCCiS70Lp24k6pn/zkp4f/79f+LevcXeD5g470IwCxn/z+TyNN2bObTNjcdUBV7ck2XL9Om7hy/WoiRZ/+4Afz/PpMeCiL49TPiHYRJcG/34eBOHx+SW5QkLFmsATLrJt/ICLqVj4MSvKVy/u2A/tkMk/ZPLrMfHU1L4vlXT96hKbrzJ+R6rZ8yzx8b5icxunYBRxTXgVN/u3tJ5MfLUfzgVUlbc1r3qFVZja8wr9kl7X66LrK72Eyz7bTPvoUuA0dZbbZffWdKABlpGgtzk8kIVFkeQ9mvGgDGutap8ew+5UzZeLCAfnkN6fbrguTkom2pJVfy+m1dSLfmN/8zSsbLv1ap+SvvgXc4z0Xfvuksf+8x/P8KHv00ey6L2vY/omzZ8+foJ8sSDjcLOFUcI4SjpspTRp4Nw1MANm7aWXKmzQwaWDSwKSBSQOTBt4jGsAL5Huew2kanNjZa319Y2F36dTSvpU3WQbrkVs7G2tGKfjZD6URZPXBTo7X7TC0s7CA4yFLP94tN+k0+Jf3BZ1CDn6Gh+Vdr8/K0V/8zbtkC6viN9JIVw5FydT10mb6oxOhX6D05Rf0vXl9XRR79y1312uPouilLodH58ZDLep0ra0dGNb2Hxz243jfzxRCIweuXbmaaZdGuGwBLLz5+qu511kXjDl89Mhw5BB1iCJbW1vhWIojf/z40eHYsSPDFRYiv8RaWq6/tY9pQlnfCIEqmqMcKuXadZ2juT6pF8fNbmfg1FmcczNGvVNBvThMAX0EU8oc5BR+RnOoD+l6PBYAprwXoIMTkTJ173TSDaZU3gBEsCmBqo996tPDT/3lnx6Onzg+/Pz/9rPDl77wuwErlOHf/PK/Gv76X//rwyGmMtqHV1kjygXU/8kv/MLwz3/pF4evfvWr0evdR48N95y4mymSb7E74UWc3I1hP9M4BS2MxthiDJTRKBtWDYseH2CNKYG4a9eugPWwjhjT4P7iX/rp4Sd/6i9k2qv6FHgQpDzOOmcm+2Ift3FKPfcOiKsAI7UeX8jCT50FlMTJb3spUytdSCmwJl0MxHt0Zj/dVMG0i5Kif9qNYy2S5QU15Z08CWtgo9PoXQp5WUZaBPy5gf/8+plzgFpMA0R2MbBteMQ2sM1dn0sBMMCYMKS+wqkbWiOMpsZSvmoCg3CIaKPAKaPPBHODzcB7lx0aMSh4Qh5ejIE9Tn493yU4Py2XLWCQdivwpVyCavvYMfJ9D981fOLpx5laSZQNtHs7AHI/0gZI8EHb3WR5NaJ9nO4Ij7ZJwa6N9e3hOgCZ68gdO35kWEFmy1cB9H0+WZcp/f3pv/LXsmmDYN77AGjvf+BedO1OhezQOG6Qoe04xdI2XG9QYE6Q9hUiz7Sphx9+sAAV+qUsymf/jXZbRD46kTFwkII3wkd1aSt1YAd0J1P6oh9sQYARetvkBDE/HQe7XQqkMDeWJsnLPta4Ff8uw5Lpl7r3+a2K0ftI0LrrtQe9NwUg5CzPed7KYYpsnLtNeXodEGnMN0+dp69WGlPqEFFaaewnjMOD9o1Us4G8q/Zwo66es7SOnZpJ/1Fw1jujj5YpfzEpvo6rz/vGeoFjkTU6t9xxw7Y19mhZmd1hGB7o3iT9FkDuks9WMiziiufX99yOkV7QLxBBqFzK0rtvZv22Ua/KGr7w8JqAsoDN/s60japjuzZCIi/t2V8ORfbeaw/X+OPMr9ria7eJSuS1tXD3yZMsrrezw7azw01pYZaqXExp0sB31cAEkH1X9UyFkwYmDUwamDQwaWDSwHtAA36O4x/6AY5DsLtzkyimNxZWVt5Y39x0Few4Sf50Kls+5HEC+mPfs6nPOlT6ddCHtj7Ox496Pu/jhMVJ9/u/+Ejtdcmwdzb/zjTPTwes6zRd8+l7z/N5fT1fzzwPU/PPPVn2a7YGD56L0RsBxpZ05ssxcrHxbR0jpxLSf6fvHVk5AvCzC/h1eDh69Gic9ouspSVQdpPIqYsAPVeJUNH5PkqE1T1M0Tx85OCwRlST0S5O8fN84PCN4QAAmg67i4rb1i3WKBOwUTbVX9EoKH3UYTu13dfuVwZaGjJSxpX/9J30oXb05Bm80oVU1f/toCJzjtnYb/llPHEWlWVJp43jwgWjcw4MVwESvvWNbw4/8dm/iOO4L3oQGJTW/l04f4lIsd8dfugHfiB87Nc3v/nN4f1PPzP8lb/2V4df+hf/cvga0WTf/4mPJ0pIwCJ6Wdocbmzdyo6DV6/tH1YAyuS7Cgim7AVYLNdi3EQ53QJQS5Qb7R49fjxtHccpdaxXxmlgDHKBnYwfcFiBH5Q7vUugZWYXqEUHmA6N4I3gQ9lsFIbdj5EdGQ/zEgk1R6PeOqmLpOjQodBrLooahyq2yU5pz4cM2QS+buHkX7iyM5y/xK6quysBmXaJONH5Dw/olEH6AsR6jGkvfJQh8Bb0kNkQC+s7pW3ApneZsrpvkQXyAXhxwatf+4iwExhQVq7dYdLdHQXRAt6OfUDZlFcfI4uIAik0NLYAQPbhDzwyPHiM6W1cK0Wmhoaqfmjf2TkTXq4dpc0JWGXtKKbcGmkqKOVzaR/dyXLt4oFh5b4TjB8gGd2Qfv/+baI47wJ4PjY88tijTNWtNea2eKaUJzvIjuuOXWWqtABswDGmUB5gTTqfwW8D4t7Ls+qzqU34rGtbjqNBY0n0URvw1t5GjylAXyNd1mWEQJDZKX7qxmmB8iw2ApZqAxryTBl3yzmiS/Ly/HHuvKap8tK1ZfOpaTq/7z3Pt+V9vUuqzebR9fo8X18am7stb5S3p0Bb1qnotFPRsHqPqAAj90zztH2/0LZFhvIpR8kpRaXUS7sAddgMm6Rm0w0X6s+UYvXNWHQ0XABO7xWeVO22nDWeLYs0/u4h8DHYt/fy6t9H1IZDj9HeH5GsP89ffViv8/1jhOXVjjpXl7x7sKemsVwJvY/8RU92jRF6WGWK+UnOJ5niu8oj1cmHsDvUedN50sA7NDABZO9QyZQxaWDSwKSBSQOTBiYNvAc1kE99HYednVs3z51/681Hn3j6FP7gOu5HdgBDJwkx8UM8X+hkOP3JpHOxD4fcD/Yx2uz2D3rrkIxU8K/s/lU9fMgrx2bPMWhHQHodRsvxEZISDIFjYDJ/3rmQn3mm5uHZ1G21U2Fel81fz/Mzf97JyV2cEOUiSomF0XcAXwSq6A7Okc7kRhxg/1YvL9cU03kWsFlhXaRDRwDKUKoLiesAbgLyCPqcfevMcIHIFKdfCqYd59A5JxhgOHb4WJzxjY2Dwy2mZgZgY+2lTSJljgK+GeVkSjTX6GzROWQsnbfcRVRO+6wE5CDr6oy6C7hB3QZWor3cV43WsaBR6bLyt/U+sQH7KYB19OjxrHcliPDGa98e/o9/9A+z498xgL6PfexjLIr+9ejl+N13CaMGFLvr2PHhoYceAhvaZiH1V1Hg0nCTfj7/7LPDH33pD4ZHH3p4eOSRR4Z77ztJG4fQ1cmMg0DGOUCLZYBFQRB1XyBK2aVA3f796P4ga4oF5HHK1dawlnFx3ahaDy5RTupR3aFHbSl2jRKcytn20v2WpnSrlspBrkgc7siSTldWeXRL2wZTaXyAaIn+Wh97LnZehdaRcpOGtCtNxrOcYA0u9o/OfT630dVLb5xi8XFAWwAbo70KGII/jQsuRY60i0BGktnPfUSHKRw/y/Z50Oi3tAuL47PE/M198Ax4Ct9iIR31IAl4ZoexpUSZpSPsTmohNLEpgVf7EHAM/t6nPuAQrD71vU8Na7TpXhP72NgSa1IzAcoabIw+eRFssH4ctTM2Pe1R2T0cf/UszatvvF5ANTZ3gMhMRTRKMzuVsh6Z0zLlKaixubnFc1nrjDnmAmU+1653573PrvRfZ9MHAbK/8JOfSZToAnqp5xSgTHTMPpGUofb7LZsAACAASURBVMdb4C3rByI1b8nkF6A2Ro+hqaYvUK3uUUvZEWOrnI7zop0YU/P37BRSExIkBcDNuBb4ogFKt2efUO6x4nIEwhhDp+/JTsDfC6ww7ZvX/I1IMxlFFdlzLQGH117SXteQv32wF5aZqryu/TmzT1+mY0uCr+rMVPIjjzYkCSk801gBW83bsjyf2Ms676brN2+xS+n6cIvluKJJxwc2joNAZdaGY5xTj2fCtqzfv08Uzj+M8BjN5LDtTYC3sj3Lqb3PKF41Bg9+NTqe/kFDWlP3gavco75c2iVp8l6lzz77/rNW1VFvIUo9NZmK2BxXqKT45bla5CW3u3iCtfhOsOELEWRlf/AponCYfkwa+M4amACy76ybqWTSwKSBSQOTBiYNTBp4b2jAr22+v5nw5fpJuKgACm/iZL3BN/W1dqpwBAgu0AuUvD7oKzKinB/z/AbXqfBTXHBr5sl4ZX5VDZ30+ej3guS19T36usv7fp5u/rrarO//+Wt5zac77y3LX/11xHCQbKemubRDWXIp9p5cXlvOmS66s93qASIe2EHPtl1If2kHB8mpa+VHqow40ktMYzPaSSd9gyiyt1mg3t0uXT/JKKfzZ88SJXaVtbZuJMrFqChBp1WBNhrbJULqIFEvt1iAfB0n/+ChA5kxV85cTQu0T/bFfpkid67m9D3TM+UKmftxcKCd12HGwL5CY363Jctup/VquVFgH//kx+jTfzH8s3/6fw2vv/768OxXvjw8961vRApBFPt1z733I39d77Co/9e+9tWAhSfuOTkcJxLpGGuX/diP/djwoQ99JABi1mQ7e47dMS8yNfUuaNeHe9iBco3pmc4mOnfhIo7wjQCPK8tEDwGW3GIKkgCkUUMCHMqpg32AAXODg+wkR16GKTqoPqpzpwouxlkuW4jw/HB6355dl6euTspWy95aH9Yxx135ehpVoq6SKwgEQIPatTnpMp0VOUyxRZ1ikvy89yyNepez9baxiy3yX3nzzLCpOILcDP22EWQ+rqLLyFegmNzg7Q95UuxzWmM6og7KIgF933WtMe1YQNtzSOS7HABtB4BA0l3Gyzakq50VaQ8mvh9abiOnXJ+t3gHQKST0Dz9wYnjqsYeH1UXAC8aKCjX1jLYELkoPJS8/uXdH17L1RE7y7ApkOY1um3CZI+xoeYkpvkZouvPpww8+FDB1FZrV5bXYgeB07AHhvXYTDYEu9XALcM3xF1S17Tx/gK/PEtn4O7/9W8Ojjzyc9QP9Q0A/n45Hng10aqLb0a/X8rDMAXb8Mr02U/IEdcyL9aWs9I6NhU1+JEJvxD9kF36ebbN0UyBN2rCA5LNvX+bt0PzIOOZbd1be19qEsmpb5tGwgFKnGX1ncG4+9U6s93fL0vJZ5rVJHp1fL0ht2mn3tKeSSNZPWyNt10mhfOiDNO/GM9LDRpgJ08Amhhk4dnNzI3pbQcHas0k9ZR1BH5FRp+TO+jWTtd4SM9m7bc/aknwKAJangClTNylTTo/mbV9yBCzu8RzHel43Csd93uPYi/ztetolvxO8VOgsA3pmhC+fxJ5P8s5Zpekk6o2kNQ5dfzpPGrhTAxNAdqdGpvtJA5MGJg1MGpg0MGngvaaB/mL2D9d8hQ+bb7755uUHH37yNJFBl/0ru8sK6dn693edP6Ntks+9U7lM+YDHG5FJ/o8f+365+1EvvX/h9rob9Nve5LmdIss7P41BPJLNaL24jW7uPo4K9/KQ5s6U9skvh0NnpaLfpBNwKL6jTDp25Ou4JV+ayGcvdeSNMMH5weFaZUH661dvQOFUGxwjopRu4fjFUdJ3AhjSkV9AXUsHXW9MoGw1EWFO3drAma8zOzZevJQIsY3jx+KEC6jpqDsNaWWJHQsPrQ377jo6rCCv/dSJcuh0RNXjdhxbgA/uTU2Tm/GHJTO3KnrCoaRPWSsObkk4cfa9oqvq2ulvRjqYGqyRfzmCAhfKuDR85jOfYUH0Tw6f//znh8997tezWYH9E7i6izW/bhHZsUIU3uuvvjacf+s0i2hvZFqmzqa6sU+Hj9w1PP7448OHP/w96cMVpqi+/OKL8Dqd3S8FJ4+hA/Xz0EMPApDdTL31m1vRpRFsTqdzDJwqd4QNENxBUF0qc47RUY39wWuZdYbMsk52baT/NeZoeMSaOsJOHVimnvMP3cuT3BxOK9WmdMAdO3Wrqh0WI/eKjhNtaDf+FDcyubOdJK3bjFXGk5a0QR1m6BYAq65tDMNLr53mmqhGAE/7QkXahkIcAF5Jti9gZksCBPATnGBEZRS+o+h1irwKDH01xoJbygUYJSjmNN+UCUZAQwRNgkrjlRvdRp/HekYG1jsCVupCvbFi3Ce+93uGu4/AimjKyM24GykVwAVJO1pR/brYutGBJmkdR58p8QHtyvHe4Lm7m0jLS5cvDK++8m2eq/U8Y8eZxnz0yPFhmQ0H+h1x4eLlbNygjo0uPHiA4Bvqmxwz1xJ0GuaLzz8/fP4//IfhAhtufIzdLgWRtKtDTLv0HeCbcUEwUkQGnck/tmXnAcA2N3gvcrnEe6LeB5wZAyJ8ys6kh+Ad9hZQxOetbAXrylion+hQ3ZOUx2HONFrOC9iwNuL7Vjm0tdipBkxyxP2HBLnXJi3Pe4MzUcThWbZik7arTdmWPxwfWxzLRj7SZQy1GwvRh3xvYS+WzcYyoVOp7Y+ipYIwmfXrvRQOVS6ARrOlM9ukzH5xSr+8INkb24m8XAs+b2CnRhR6llb+LOVojBebq2C/nLUdx8Vy63qG03hw7eClL9VneURO6PKeoI73CmB9+xEZGD+jpU0p9zmjLNrnOfWPHum8TZGqXS5af9SNPGOZ09fVu+PdclpH8ZCDYsr5tcSTcveFC+fu3rm1kZ1GIou9wGi6nu1NadLAu2lgAsjeTStT3qSBSQOTBiYNTBqYNPBe1EA8giWmI/32f/j37Oz3xDmQn7M4e/nTM1NuxAHyKb/slCs+0suRwckQ9RmdOL7RSToQfJFDp6vBl3/os/A41+MHuyWzD/3O6w/4ONPQzifz8hf1sZ5lOghdt2nvvO/8Pnd5gCUFhkfAvxmvcuws7zY9myKfjjB9XGHtIB2gJUBCnb+AgIIisNzG0daRkYfO9iLXukamAmgAz/athv8BACEjybKQP9FUrokkUORi4zOniXquhaWedYAX8YqWuS/wxYEpx670oVMmCFhOXzlnpSv7oRzRQcRxwEouy6zfOm09Wd/rPUqqkJre6+hlrBvb4Nrpln/pp/8yO0j+GOuSnR8EuNgDgo0HriZy5/Tp04CvW5kC98pLLw9f+/o3hjfefGt4nh0w7yI6bD8bHjz+xJPDM898cLibKDHluuf+ewKKGOHl9MrTp94alrFZZTE6TxBuEf0YZXbo0BEW4D8aOdYAMB1Bd6J0nSUdW3UJy9S1vg549b10gOnbtdiyTvliprOWw5sC3evYffWfm5keUi4IZQPvSOiT7AI0sAuuBQCETVIAva0kAsu6OMzNJ3qmQsaGfEEN1h4fzl26yswqgBEdaOvYW8GwAGEyTwMVCcZljV2hcfUcU8WK0OnAK1RAOB9kEzasOgSjojO8KNckc2H5iiAzAwKarA5RD/YChFGR9m+nqRzZAclWl3eHp554KNMrXb9ukzFN5B5jI3AxiyALS5+lBaKBNoZtpspZdvTwEZ4BpuICjB5YZKMLQNAFNm/wvbO4+OSwS6TZ+fNnYxOPPPjQcP7cxeE4wNYCQJWRhZfYJVbFO6251FRgifIJpB0EADsHGPsbv/qrgG0vZ4qvU3ad6nuc6dLKYEp/OC/AxGdL3ZpnXzLtbaTJc0i/gcpT7vswdaMgBiXJZ23vOTRLGo+eSpmxjYVUDcv6me1n3ZIa473nuaj3fnbgke8w64c/YjQvRqvSaOPma5/aKU3OypCOOgJQJWdPG5ZEGeZlEmALH0bYiEPt3mQfskB/eCkzeVWUn/1stmy+V+9c06z1pD1rw6zFNdy8sTHbudK6Xd/nPzbme4DkSPZ4el8yaqve1HPu2PYfeZqmeXpvXz26zH77HpfGP6KYlFGamf7GPMtaNusVn9JVxskKPEutS8/ysrr/qUvWDhvRAsPvWzz2+PseO/69n/r0/j/+g9+jzGc49ODSs1G17pQmDbxDAxNA9g6VTBmTBiYNTBqYNDBpYNLAe0UD9cmuMzEmLrZY2+of/oP/cfj1X/t3V3/253/hzOrBI+f5WD+5u72LR4EDxMFHNrtZVhxRIhlwDAVqnH7mNKdK5Vj7EW/UTj7R+ZO+oI0+hB/4fqx7SOPZ5HXfezaVU265tPHAQ2OZfEx7tPCcdayc1abptc/a8Z45M/RJ+f2XNDLQgaoojHJ6qnDvpwEZ6bd9h2QZPluwcEqdkSW4RoBkrlXDVDUAsxWmSppc40gHzeMgEWFb6KcAGBZcZ8rXtlPb1AOOzQbTBjMVkO4vMaWypvhVfwPIqUN4AkGGd+tOVMIcx0ugwlTRcgJBpXsyki9dxqGGIG1b0GOypyf0GR0ZJVGp5CRCxFsce51jo4O83wbsEyBxB8lHH350WHys+qx6ree4CFQ41fTUqVNE6rzEVMuvDc+y7tjrp97MtNOvMD3z3//GsaxPdv/9D2Z6m1PbrG9kyjJTJTWdZaKHbOfk3ScypdKokIMHDwfErOlUhFYAcAmOlLONEyoQwb8ed3x8QE60k6nG9H/03hsEa8B07HnprPusLjHsGgv04bWOKdnRowrhRl16b9+d3poxMd9OhASbG3XT45KxkX/0ap3iuY/1vlx77cK5q0wTZIovcTG7gIMYEB3BWRfI1ki1AfkHDDDicQUbVUY1QVFCRG287Vy5lQfNIG+PVR4LnmHH1BgckyBwmAiikK0ud4nqYo4nN/AwcgdkTa2nHeRw3TLfCPfedWR4+n0PJ2pOu5fcXUntr/IlKos2UDHgxeKweZMps0xNVnergNNGGvr+uXLlGgvdA4wBlq2tGlVGdKXl2MQbb7wxnD1zfnjz1OvDKut5ubHGMda+E/w6zu6oW0wJFlSlQdoHvKL9RSLT3Ln0leeeG375X/3L4a3X3hjuv/++4SMf+cjwye//dGyR3oxqtd/1/hJAqVTPXsZd+Sn3EPD0HHDGPNoycZl8FJSoIs3OPjcglghOx8+nDyXRYq5H/JZr9AuT2JTMRopZffLKhqzHkGTH2wLPA75gB0azyafoPDuSleRr8r1ZfbG9UeaRyvUSu7/ZrVh5lNVnQBskua6Z9/Jw3KxqnRz0jd8qUFkmta0rUyXvXPNRGxR0Uke9wylQWepoY7Fh+CzwrN9iSuVVonrdTdh3/wr27ztT86UneRZ9AhwPk3JFAtp3aIxAS9+VkfLqH5XpV65h5NTe0oljCxF58lZXt9Cp7wzfxfV7q9qwLftYXJnmq63ToLbfuq62il7+naTbG2flpLWS0x2mgcjQMSI89fQzR/6fX/xXB37pF//v4e/9V3/XxmiTOM/o3t5MadLAu2tgAsjeXS9T7qSBSQOTBiYNTBqYNPDe1EC+nPnsH155+YWbly9dPHP/oaNEke07ynf3ih/0+Eq7bCXP97szOsrhC0jGdZzG8dt7r4w6cXb2PvaNrppPfvDrEFjHD36T587z3jI8ba7KOfG+HQXp5mn7unnN37+TVqBA54G/8tsQyWgyU9rk7J3lLVPzSx0q6xAKfm0REeNOfubbZwGS7pt5OnZxmHCivMdbDE8dNMGd5WUdKndfBFhKuVESpRvzBNb2L6yWk6cjho7idCsfdDOd4Dlbv+VvPXlvfiKT5D/2y+HpvjVNCvnRPL1vfu4EN5/23LfRYRvbCS+AB1diVwaruSC6GGf6BxPzDx86Orz/qaPDB97/zPCTf/6zrB91HlDjzPDqq68MZ12Xjd0+E3l25XJ0cx1Aw+l0hwEMBUmOMhU1u4ESUWSEj2U6wu342l/7l2lsyobelS3yqadSRQCL6Ar6pDHfunWv/Xd0R+lDNcJq1HeRtZ7qbi/PiJcalz1dplQ7ACRFeykXYDXJO+MVfTG+YNQz3jbKsUSk01vnLg03iKrat7ifPIhl5TkH1/LDxlJXsJr7AvC649CaRptIOJW3AY1GkCDF0KsbfH5rLmDzOwBWTruEiv/qEnsV4PX5bXwDvj3eggegBwDGt4YnHrx3OHFUxvDiEBj02nYbKIvMoCL0jk0IAI85F5hMtBd98d7Iyw2AVqMLZeT4C6LGNpha+eB9l4e3L10ZdpjWe5SoRqe2HTiwFhBsB0BNsE17yRTojPXC8Obrr7GL6j8fTr326nA3U4IffPD+4ROf+NjwxKOPpX2kSJ+UT114znRTrtW/Gul8KQy/NQLRdqRNv8Z6dlsbDGDmeTTI8O4xGWn3OJMxpnlebV+t73ke5pVlVUVBMIEjx1MwTbNJ/brizncPsvbzMNeefFtOO2y91B37JpCljkx7XbAF22LU7DT2kuTzyb9txj2AHZnyqr90KJf8kVM5xnZSM7fYHPndtjRWlfXmLXYmHQFVaaILOrvIrqsFYvkeYFw43FAl74ixX2neH1CqIJ+ZgP+WM5625/vF/E6lE+2g+mm+73zz5e0fUzqFVk7w8do0z8v76B5e0cVY3rSezU+dKEO7kU/xWt/cOrKztXPsM5/5qWHtyLFh/eplUVuq7MlrG1OaNHCnBiaA7E6NTPeTBiYNTBqYNDBpYNLAe0YD43d193e85SuanK3N9Vub65sXAKXOEwH2KKDIyvihzkkKP8Tr4z47Uw61W5eOgCDQIs68dH0kiID7RIboPHvNoSNs0mHJR79ONo5vtZGiGXijF6mT0lM1q7R+tuPgnbzcdY8/qaewnQk7Vk6s/C0qsKPdRkSODOOyavHPBFN0eHREKqJIZ6c8fx0YnaRFonU2Af3KLyoHJBESRAa4ptEtDh1jz8qiOyi/HeRzvR8jxBTVdXGWiHJZHvtvBIMO1hL3OnKJslkv/SyODp185Gm/BICcqiYQY19b91FCHL3qXwE15Ug5jjpNMx2plZGnfSg9lR7vHBMIU2+HkIX0DxDP8e/6titfQ4RUN9RmeTFLsTYKrePIWf/EiRPDyZMnh6efeSb5RiVaLnCiPozakM5YOJPRQrbjWNRZfanLsiNlM5mXf0Y7jU610VCz/mO30lTUIGfpSI6zfTdipXUaulJO8up+dPxTa++HddI2Y5gUm5Jn3TK82LU6qgxpTdk5j+uKLnN8x/YdDsZ6AWDqFlUuXr7Oc4UOjBiTKXSmjJdGKVqRcabMMRv5hGjux+y5Uwx1JZ3joh60qWSbPz7b5NXOlUjuGPMA4ZSPOhRFq34U8AMobvk2C6ax3tywcW34vg8/yU6s4GU3irf8fXaN/qFB+O1NKzTKRlEy7sh1AEA5dgata9BdZKH9xUsXh7WDB3jua7zUo8DpEhsOHGHHV7ViZI82l/Hkej9Tbw9TR16+t65duTqceuP14bd/87eGdaYCP/rE48OTTz45fOYnfoK18D6MdETgjbp03Bwq5TLJQ/lqmMdM8t0R034tAZAE0B51W9qpPlMcvSkbVOHXf3jITX4UT5/f2Bt58tVu2sYkq2vPqZR78wQg+9ybUPhHh+SlHjJQx2Gzqry98pnpZP9Gcwph2WqNeWghVcrwpM2Sr+7DXLvlX7VZ/bRGNnBgPNSnuQZe5Sb9s3XHTe2YDQd4z4A7KjkdWjlj/5y3eHleZzqu71wBX8fNM+JnjOyH7cY2ufKZN7nOFwt1eYWM1e+Z3WWgpZOPZbarzIJstoFl+EccitSL9iBIbQRqyV38qMgj5XgUXezF8bEgSf3s8bDFjDeZ4TneuwutiT+r5OyfraTTjleXFg8COB5//rkX9i8vr95c37dAZ200pNOPSQPfUQMTQPYdVTMVTBqYNDBpYNLApIFJA+8xDfjpPPf5rCc7nMO5PIfruwH4cGiTKBX9I4EiwRgdhQKCqlqcjt29be29d+2VMNah8R8f8DpHJsuNRtJVmW+5y5u2nQLJkhdHpa7Ne7cUWeYKmtdc1kyWmaNFYbftOQuYc+6/upuXozxgruXGekU46VvqA6BmG4BgiymVJmWQvtueOdDUN8/phZBk2p8AogCP9DPZcdrCAyfPfJOLlOsA7e4ynY68RaKz4uoxTU64yLz5Q6dNF6rTfJm8lakjMKSxXNn6umTZGzPznVw7D1RK3327s77gYwOMMJ7xzYU/lJd/8rDY+k7DdQqVYGGcWNZq04Fu4EogJyCsOy0CLNm29Rogg8vIr0CzLus2vQedRfE4uKXW1O+Fx+UTvYzyzsutnKkPs74u2atvrYduy7PlnSLLaBfdttBYU+g0z8Zlrh656KBBp3qOlIuAvOHbr78BB8Ax+rRjlIpGpYMfJ55LzgJZ2UmT64rUqo5HtkRmorXZVMuStvvpXfcheepvzBPu2MX3DgghKE1+aHxGY1s1hpa7DBNQJ/nsFMlS4t/34fezc6VPUEWUWkXUwA0KxiYCSgvA3oK3i60L7Ow/wLRkgFLBHaeuHT9+PBFkFy6A5wOSHWFNsdW1Zda2Oxi5nT6YyC3BEvXCvTpue3E6rnZ69vTZ4ZWXXhyef/Y5pmCuDj/4Iz+cSLRPfupTRJA9GP1kuvNsXOpZa7uBOXL7bBaAMovUFNBarOe6bSVnpYnOC9i1fperw9Z5nzuv76UfMZwZbT2vypGRkCTJOgUeVZl6ExOSzkOLSZ2gNjW+Y9VZ/ebd7fe9I2jq/L72NRlwWfu2/QxwSPPDvJKzbN7xlKYAwKqr3atTn5Gmbf7ey6P55J5x3R75XGUNxw3WoRPglUcB6fLjnYQ9Ov4eKMZmwqf6JN+8TWdtyrvaK/m7Xe98H1rP95b5SA4tVk0Em++pjkxMHZvi6PrdB8/y8Gyy3Os8EmPbAozz9FvYc2w4z0t+L+wrm1aPYMgr++87f/bcPQC0r/Ny0PhroOpcDaW16cekgT0NTADZni6mq0kDkwYmDUwamDQwaeA9owHdIZOf37PUvlacRXI3+WA/zzpG53dYQV4wJ9FMS4v4lziYEOhwx7Pgzt3/bvGBX04A3944HdIt4ayQWY7u+PFfq5fpHFbkgVEqBbiM9WcijU4b9+1QWKSgcShGRyN5c46F9w1UtKNhnin18FA868jqz9SBjGN5LkIttITjAq18TNbTn+p7nRod7E2mb4m5GE22j7Cecg4LtNnGmVcXysQpYAJ/1R8jUSouwmWvDHRKdBwk8ncqWORncfK0HnkLvIn8ATsAHZjWKS5innQCSOEDsBCQj0wBOIorwdt/tT7QmGe9uT7Ky3WFlJmaVUbH20gcw7Q3nuXS917Lq9cbsu9GWagT81WBZyPBrINbaBV4K/1om3jvdF/C0AKvDEurFR2xt+6P9Sp6LU4vnUxbKMMIQlPuQWY8r7BTYfo1OqLuxBgH2WZJltU5p1l/BFgcZ5NyS7dHq27K3pTdaEruQtv0fWPdTl4LAprEl7wOb3RROq/7ooAWWS3f50Bbl4Il1h+7dv3m8NZbZ1Jf/flMBqbqAdeGAMdSjzrhHQ+o+lNRMo4ISf4c9q3OYz8cd4ulse/YnWeTduRl8TEjVJzhH5ujUL404fvDZ2lna3146gOPDE8/fmhYBnR3huaexsQuBTTIE/CD/y3ONzYKJA7QpYz0XdP0vbHI+mNX9l+B5sZw9vy54dy5c+iGtcgY76PsXOpaY4fZOdZoIcHstcOsXUabrl129eomUWSrsc01+AiEPfDAA4nWNPrsoYceYk07FvbHeJfVqdF06aa6LpBaYFF9oQXO6Nsu+94be1VTe0vf1jWlDvJoVj4b2m+vU9X6p4T8srW2vy6r/FSOTBl7+Dq+o4SRQ7BJHSqf16YqR8cYnXxMfU4/4DH2hnrYJ0IKMGnfluefZzuauvZB/sW5XxKyjrwjgDOWYhb+3qDQRkw2YqKCV/LSnmLHZpNpJK/yqsWQc78AiKUE5vMqQTwlExzaHa6xe2k2dPCFS75r9Sm/z3tFEdtcye/7mzuOSmkbHtHFmF/9KADLSFJ14nsrsiq0baMPZat69e4JqM+afKmj5oKK741rtxE+yFPPUY25+trLJ483p/cBOqF1M5KAvfCF/z70v+B7ToB5a4G9L/YtPvDAQw8+cPXtS+cZ9escdjIq5rzXYW6mNGmgNTABZK2J6TxpYNLApIFJA5MGJg281zVwxwfzzjrOxGk+uN/COdjQQdC54MT3OS7L3BRKgRyWTZ45Bq3IgA99M3eOsxEnqJr0i71474kgTadyIvquznEY+d6fpytHrvLiSOjoxZvaq9v3nl3zRqemHSbzUo5AM2dvrOq9kVCWC+jZbsmcqLpcD6yrZJ76INZlJpt1Ux+nKnyp60L87kZp1IGOmwELARCgMeksF8iFY46z77VOoE6+dDpCylDRFmpw7Hf8n3L+VKE0/ku7tqP8Fswly9Jv8ubPd9JZRZ+4Hddm0X3re+s1n7ou2ZSx27+NZnRGzXOqlPpNfzknIbNpi3L7Hd44gS239ZBs7GPJ2D2UtmWpumpjdHRjz+XUljyle6c2xr5o9jY5aef2NktfPRWy2+k68/fmydO8OPvcNyBS3WuJtQZ1XLzDi6LIQ55JHtaFw3CZKJkr19i5c+kITjE6CIUVtKtKLUfWm4qpUO555i835e1nba3ltt+RZczTDiIHVbwWn0g79k9jFkiqjqHEksoZXmwtmeMnfvT7WTTfukQHYc+CkPJndEf9IB5524AftzgE6C33WXAX3S0Awy2iNTEIaiwMdx07zrS6bXaDvTW8efrUcOntM8Mma/Y9/ugjw1GmUO5fPpYosv2sPbZ/ZTULo68Cmriunyk2PKxkuqZtmdw5NVM080wja41K+mVfow/HAp2YzMsY201k7dT5liV6iB/CKwUwlW13fc/WFZDqeq37bq9padlL9F2y5I8MtNGywZrs7QAAIABJREFUNX2myYZy70e1Md7TXsxirzhX8oE7R70fvN879vonsfw67bVvfWUr25nRlNghTxvypXpZSfd/j6dPrGl8OqGFJ/fyC1hEnwVOt/r3AZGlN66v5z1Zz0G/f2uTFKMA3TjGd7VjMnveR562ZZJ/VNCScd+/Kyy3rjQZ8yI0e9T/CJCN5Rn7jI085xQAfbWjbn1mHfvqr3T9vpGvumzd9jm/I6Dn3UZWUupAvLZvcemhK1euPIT+n0e7AGRJpcbxZjpNGrhTAxNAdqdGpvtJA5MGJg1MGpg0MGngPaCBdkVu7yqf5X6Z882tU6N/uX6WaSlnr63fxGNkDSycUj70WdpLAv5qzeFfxHdwcHVv4sj513zYi6G5ZtbSEguHxxmUp3RQzgEfOgM2al6vGdUOgrTKcruTYN44lUWvilTRDcUjsrdDg0Nh3XZk7uSLvwIvnZyi4SL8Zo6Idccseju2NWYARnSyzSWiBHbZEU+eRpHh9cN7dHZ03ADjttWXIBs60jlrl0+58O2RFR1vrEOjy180AgKmRRzAJUJtBMeUwKmW6Zt8jD6RSF16IQHyCTd4L7dOrQPPHu3ceX2nrt9BW600q9A3D8/No/lI6HVPOVNeU0XLIBi3cTjRV9pCL5m+C02Neek6TrD1RrMNf/Sp7KaibedRO+TavkXHBjLV2OET0w4HTaM9NZxxMJon00DNi7zYDRRqkFvq2IeSxfb6er6/1tsrUy7vR1CJsi4vW+x2ilfWOhvbqOmuld91CkhBljFiKfbpNceFt4mcYrfQbaYshl557XcJnrwFIsiwhGEfNoNWICi9ReBZn6t/AVNit5SOfW79BrikX9oqDz42rQ1i546rh88ESt7HVq7q2F00eTlkGuUu7w75LTGI9508PHzmBz8xOIl70XwO+Rj0V1oTXJCn9gw4xrMUG+B+iTa0fd4AkWEHIE6wyTXJjh9jV0qeD5+Z+zc2Aqrdd8+J4bEHHhqOsTh/Eg/0CuX797GTJzugrrPJwS2ANhf6t02BlqMs7H/k8OEs9u94OTXUsRZU6TFpG3YapfaW5yjjzdjG0OgbXUDhaj718p4hKrPGSVsvkarX3XPzaiwdpZr2Ws9Hty2FY7LLOJmXf56RNXqas1XpHJoyB9uQZ4GRsYVkOPYld2SUmOTjpe17W8+a1x5ju1xn7bDx/SJt2sPaYjOjnWnf1uvnEHVFoDy+CkcPtC3bYYhDu2XEWolBWbWXsVaf9E9+PqOuY6n95Zn03crvBu3jJuPPQvUZC4djhcZcjL+AyYrONd/3RKZIKh/RmeET8aovtJa2jCA0TNN/vjt8f+eOer0WWPpD3U7hhX2U7qpf8kv/OS9Et7ZZfVL3pvRNfYyMMr1cIpIgv0meAntZZ9NnAENcpv/ma6ekNS7v//0v/d7925sba2bAWJ4EcY7Mkjn9mDRwuwYmgOx2fUx3kwYmDUwamDQwaWDSwHtXA/UFXh/Qfpvj42xf5GP9PH9wv7mL06FrwOc9vgx/w8dhWFpyyhrOiY4x3/b9F3k+46NFy03z3+NeO91EB6qTDsE8Td/3ed7BkK7r6rNY1nTy85qf4VfX6Ujype12PHe92kGwpDEvznnd8nOsM/oUARqUl5IZDx15yuOccO0ueq6ZZJSYSZ4B9dK+snVEg06hUXkli85PRa+UftwZMzxxxgpsrE9X89RBHbp8lZzeJ1gYWXCWTNXHKr/zp2WmPve19e9M4aP3Suo126Rr2ZWl+fR16ox9a7quo630lC/zwle9jjxrrEYbQczk074ARvP33PX6bJv2fD6qx7otS9HZHm3BTx4BftCp3mPLIt186r6Z19ctx7vdF5/b200fRllKdhrUgeZfort0kHe0ZxpBROkzHZmzKbJSaLk5WwAQr7Nu1o5jDVgmYJCxkcBn0mNM32197tv6HOZ7erWs+5eIMnTW9hfulIdGUC6gMMBCosdKfnULQY6A6Tvrww994qPDY/ch2A10KahC+Q5ne7UNf5+DAiUp85lgTb+WwzdQXyuq0x4F4qx+/BA7VHJ/dP3IDEg4cugg64kdYHlA9INcgmfqUUBO2NT7jc3r6aP9WgHoFhxbW1uBdwEO9t82NRFTXY833AcssYvjdQO60sZGqCgPIRXbMKUPnPs+mWPf6lqaeo92++b3dT0/NU6tD88eJs+2JIV1TF3eNJ0/UqXcvMAoqdHy7dlDyosdY1ZTS22yeFclr8O7RBk57ZUh0diPAoHQToCeqqddj4DXXM3YPnzViP0qEW7vl8Ck7d5iuvuNmxt5HpzSO6PmUvDIv1/4+8vo3da/9bS7yE2N0lG0B7H2Ijhb7+PmB1lS0Vqncxx3oh/h5+L9sQ/4p3+Rfq9e9bnta68/LYcAnrbtvbTK27pQDq9d55MzUvLnl7GcFgTF7v/Yxz/x4JPPfM+BF7/5Jwgoj+1qZE/U6WrSwG0amACy29Qx3UwamDQwaWDSwKSBSQOTBvwWT4zAcHP9+s7K0sJVnGtc2dFpIGpkt7zwfJz7kZ6Pd8r9OMfnwDEhgkCnXweBv8rXWj3l2vCdn7/6O6eQT/2ou9broR68dVq2x+lFDfZUFEM5CFawvZwBAAQ5kCzOp+CVbaYMGnA8XU5wgqJvR8byvo7sOB6e+9qytImEiWywnfSqnNvSTgFn0rVjZf9dTtp1jpzGlSlgTNcSIzBt47gZzaNTYx3ppdUhNYJpl74rgw6eVRZwsm4SlSbwsba2NmvH+okkA7RcYJ6aO2UarFGOuU79CPzQD5NRa7qVc87TrK/yKppytqSZT8pjir7qMvq0nnnSe9YJLId+T5fW6/qeHV/Pe3KMDEdeDQgI7ATs6fqQWU/n1narre7bnv63iaQKb7ogZ3f0NO0TeIJ8l/qRGR8xOhn5CvzIX1vplPvYI3X8N9Nl6an7Ib02YGr5pE39RNBYVjbZukJrDEeNtf0JOAaVdRC2+qg9wCfNjmLlnp4FTKL+BvK98dZZ1uBiEwOmleHGxxbIUBwZRh8CyfL2sS0gruQtkr3nCibQ0abPlG2PtrCLPclD9Rj9Ik0U7BRHZSYJwGXnWHWdfvSzSSFglClT2Qgb+5t/4z9h/pdAyFYA4S0iTQ0fq/6qXxZANLKMpLxGBLkbYQBg2rEvPuuuPeYYe9825U6RRw4eipw7LOrvYv2rRrKRVnjWUF7aWV+vaZTWFXQ9cIAxoc+HDxzkei025nvDciohkzqo++hDPVBisVFklWpNsjxBFLgBSYMjlmtz9lFYSODTWt7L33a8rHPJGDuxYmhoB3vyGfE53+PLc+24hyzCoG4BRrl2m7EM+NRYV58sK1vre9f0qlo2OYI7sVPz7ac/S/+5cpq9+vRGmyY5xt2OHbR/WSsMuq6rxOm7Fej3QmzGuo43/KWlr8Wx8uxQr2lovwQbTdIYZVjX2hy4K7tX3uRdYDSj/Bx37cPDvuaaLjlu+R3k7yzgJafGR154S5c1GpUH5kbw2lZs33JE9HmSXl1JP/97KuNK2V6bETE/GkBV7Oie/jqe2lj42TbKqPaqb3u17RZrj8F7VAGnTBlFgETuMQD0FbPmd8Q9f/7Pf/bez372pw79nz//vw//w9/7b2CjsWYw5llO15MGZhqYALKZKqaLSQOTBiYNTBqYNDBpYNJAaYCPbz6iy3kicuk6H/lXdWnyUc4Xtg6BJN7rAMRJ4ru7o3bkMtKWA8B9ORDFv651mPZS0+ds6zoeozOW67GtvRrjlf4D3/txOpRBr4PkOQ4O1827y0Iwl98O7u105aToT5ifureJXG6avOLc4I5GF4mqwBnHKWcbsTg6ro2kw6Pj0ryMkliCbyf566i7YPT65o3Q3wQAAVEbljgbQWaUkIE6WZSa9gTZZGtEXmSHp3xyXWpIm7ZravAwN+OPlsdzyV9OmsVd1vSW24/qC1y5N7Ve5+m9nk91PxNqvih84hCO/GE4Kw/P0ROctwcJuo0eP+1PmQRPWg8tW9/PGM/Vt7XwGpttPaQOeVjVrK3mJ59u3+vmb571vW89WW5qes+Wb8cmyLcNx83xJhUv7WUUKLno2+ljSmNdnOINNoN46+xFnrvFbHhAAyMlJ/1g6Expj/uCnOo5ncmiDNJFFgEP7zUyQC35WRZ5GXvRB64DSCQPmdNCAQxGiO1uQiOP8NMe6avOP2DVAiv1P/m+R4anHifC8uqtYYvpxAK9HkkIKBAmsCwIqIxuyNDAiDSxP2RaCuhRrlwBFAIhROsAmoGn0S7gx/6VTMn0uuv6HPVz0OPglEvldJqmQLTT6doG6DBVBWeBZLg0hqnL2u7odvGnmW7LNlrH5kWe0T4FVpTIQxqP5tkydV0ZW7fprNRtdPRpysILfiP2IT91lbI0JKeuO77PxvvmF4LkKQ9/wBjlZgDSfxpukpxn9cY+cLot2bY0Ted9p5Rpo/BOuWfeaU6XDBiJDfJrJim7t0LrHxHUq1FZWFhFV3KWq7rQbgVwr1y7yqYp25k6K++8W3gfO4bWVTe8MVN/nI4YGe6UTzpTy5+buXvp5+t0uefSPRuDsM7dDFSb0998PfVcNlntWXc+zdOa3/eeC1ircTYyzmIOtbkIm8OAyyc3tjcPfPzjnya7xmJuGKSf0qSB2zQwAWS3qWO6mTQwaWDSwKSBSQOTBiYNqAG/tJm+9frrfuiv48BewfndAsDxr9L4CzWVgy91v9bj4PuxrpOywBo7CwsV7XEL53aBKWNLY2SKERT98V8OHK3Ign86CX7Zm2qHxNE74l4Ho/m3czDvtORaZ2v88vc+9BGPH9w3ffEZHT0d1ThB1bJldaTKXL9wYChzzRidDKNaig9OGanwxHKi2fCTKZb7M83SKT9GsS2ydtj16zeih3UiGwpcJIIGP8jpY2tEAAmOmQQIvN4AUDDizEXEnQ62u7AW3S0nWgCghIibDZzAQ9RRlxUlNTrF5SghqUAHBBkb9WMLJPrdfa1xeKdD1vqqCrIowNR7r0130sRJTX7RtIMpgJHGGQfP7mhoElBJ+0i6NEbWZexw76Lf0UHVZrqtaltbqzGdz19wDSHq2v1dQRY8RiOMtK20Z5teEy1S8pihM1v8QkO57SkXy8AnashnwR7L505Z5CetckVm+ZP6us59b5TdXFuhlBiJaaCnG+ahSNk4LrKExrZ3jR5B6AWm377xxsXhwtWbRBHexUhjl7duH0caS3s500fHPVEv2FiS0UGRnQFBbv9laP0x9oNGaZt81UYrWSdpLE+0kOXwNbop6AT1Ennm2ClvIsMAg1epe/PG8Od+6FNaJeAYABnAmIvqB/xVIN4T6ocqPGO1CL89ikzKZlu8Q5bth/KMz6EEiSjiWXMtQNf+0hbKNuQgD/rEpVMwnbo8H7W3TB0jzwKCwYP/kdv6Tl8zxSZ4nuGQ+7RfrNNtM5XBOreQPfYzgmRY4gjMUI7Ny98ORCbrAdz0tXza/vJeyX1FKGXqKve2oSrSIX7KTh3U2HDpe1awPNnkazG2JwDFGQ5pTxm9zzvY+spGXfmmjTxJyod9+8wY1eW4qkiSkb8CUhpHgUCRJGXS5J3uGEEuv6axX96nz7arfLJxjMa0HbB4bEfalFuvbFApuj8Cx4KwctkCHb3KphXaldN13dBhSWCMI32N/DYCB4167KNt00xk6D/0SG9Sr+m3Nk4roUVXrj3ntWVVf+zT+H71Pe4UXstyKGE1kv62DnxjVder/2g17bpmpQX+S6J966DR3CYyz4q0p1FtR74ItrNnU/uOYAwHLl+8BI06Mvmz2sjt9GPSwJwGtPIpTRqYNDBpYNLApIFJA5MGJg3coYF9gAtf/tLvD88/940bO9u3XIvsso4dzoB/mc528nz047OWM5UPd7/T+YD30Pktx6GcDB0RaTt5HadhdCaMAMs95y5rwKUApXI+5G1qGq+7ntemvpc2jk1l3/bTMunmZTLv3fgLjs2n4l9yeG3SWdPRtP6NGzcSEeBaZEcOHRgOcxw9eiSy6KDrNEln260S5fRosEy+0qhHr51mpg51HG8BjAms3SQCx2ip7mN0qCxz8jYfZTR1WZ/N6z6bN09vfudJZ+p6tjlfNs9DOsuVfV6/5knX5wARY5sd1WOZqR3aXONOqttub16ulkc6r+Pfcy2Nk3jl1w5ly9i00ivfnfned77Xaj5n+XPfqa+7j/P3LVfndX/6vnlEZnia7xEwj3ZMt9HynLjWWOftYEenzl0CBHQ6JWOhIQmCWXes73leNutGrqbhPJMzLjs8oEnojrz6kA7+BVAhJ/mOR9pBrrjsY1vZiKONeuyDmyUIjqyCLX3sQ88Mt5iwLYApiCEQbMTYJguqe23kj1Fj2nit4+czMr4rlHvk2Xrw3j44zm1XgmMm7Ss2JkgXoE77EEQDZOP9tp91xlZXiNoUIEOfRo6JgTUfaUs/8h95OkZc239l6MM6ptZny9x5Wbg/wGzISrbwqueocotnX8/qOiZzqYGzbqtAoxpr8zp//qw88zrzumkFuTyavvvffZqv1zQtjvfqovNLH+/+nHQdz00vuKNsPqMVmfxO+avM/vkuBHwcGVVbNQaVtTCsu/4Y09IFCS3PAvyMjeO6jB0uYxuU5P1i/3KUWc1kulNX889ut6n83+2Qh1M2pde25uuN4u+1R4a/GVsnzVe6zuv68jX1vWdpWmau8zvZe383cHuIqMi7r1+7sbxEdDIZMigm4TT9mDRwuwamCLLb9THdTRqYNDBpYNLApIFJA5MG1ABf3NvDv/03vzh8/U/+ZONnfu4XLh04cvwSH+PHcGyXXJR/1/VnIPQD3c9tnTT8j9q5jnwdDz/c6yw9RNTLB70hImNdP+QrYqycqgA+emt++BPYEh54N/twLgNUyXOs285BrXGGNDr0pvJecehHR00njHpOr5Gfh3UXWbdpL6rBujri5XBIgxByg125ZN2ePor90WErJ4t+IbMyGnFy+cr1Ye3A/oEJXpkyqXcmXFOBOzezvlIcN2NOkMPDpCO1s1ALict3a1yHyQ0StpkatkXeEo69Ossi44sbARG2dPqQ1zoVGUNb0OD+kbfXnwRMOFxEtqRNMoyeireuACEonecWfYQn9J7bgXUtKGUwr88ZJ9uHtpOOZSX7t+fE2V66jB6tn2ARbWMcv5K5bCT10Z98mSQVm0OQApJSyHhSL9NMUfBoHbEfecvcMdaulrBR8wQ+TLPIMoSp8bba/DXtaSsSc24ab2vMWsayj9BS37E22WrO1I0suuaU2xd112nG16Gg3E5m90LkTX0tnrEpW7UYfWBvr775FgvMAyQtMg3RNqXXVtHDggt3w8qIsWqbfo32XExpRIOMHNRRVySoo0/7WxnKQ81R3oBk0QV9c6xTxilhX/Doep4Zl/SNa6O2Th44NDxw8sBw4xqaubE+uDnuJjx8dvY2xqh2fdbVRcle1+5g2frz7FTP/5+9N4nVLUvTs/bpm3vj3mgyIpvKynSVq5BcxsI2FJRLJSGVMU2VEJI9gYGNPGPCBIkBAywhwLLExJYHSDBAQozoJITsQUl4AFUIF4XBTTXOwpkZERkZzb0Rtz39/5/D+7zfevde548bdlbJDBxnrXv3Xt3Xr7X32d/3r702/Xz9lqAY853EyiH4sgfYruaO90H0nPNI+j6wpyCZxwuaYrmjObGj6482r6QSHeJZzJHPzRPBl5QaV5H0dAJPjcjFPE4Q8Vp1zG47WDqd1C+iatOsLELG832m0Sj40jfchGQK1t2I3AdKJzNxf81f8P0qomxQ165k0r/IQVtW0aEoVGpOFh6MmG+RL7x7uQhckWgrfTWONHjeLtcoUIwTr0gmmY7wyJnl2IL7AHDwdDAMeJX7vw/mhU2dGEOxw5aqM4NPXp55g35WX4m6kPW6u4KgrObCbtDf2+e+CF7Jzv2GOeDQmWA0DZzCi75KJRu3Sf5OsEovtk0OD08KjQV/C+DjgGbjbToaM8uChFKAvxsk8rJHCeAv8YKHEpLBfbqnxu65H/DXZYu/ZcwnvZus/dKECl3b6Vj3m6/r+viaVP9ASmsJ861JM2tnIcbpzltAU3akYYFhgWGBYYFhgWGBYYFhgc4CPDDzM7Qeu1fTD9773sVHH37wqdo+03FJ0ANnQI6G4cDjQbw9jM/lcnTKASiYeujnwZ2DlGBKj6+QkWls64GfROANWhw4DEmhAS59JMrl5BVUZKpaOV9pg3dPIzDkwAQu7cBGp/Qlp51FK3mti9ciX758afrIs6fX4lhNdnR8UF/Hs9PenCDxgnZkgR9l8Fh1Qo6silf6VTRWkFFnddap+JBHjji8oUV7aAcG+n07dVL6g1utJUvgcZJ7epTp89h0ObihswkfuuFnPYXbp9CljX7qgcsYBL6HhWbRLeccqn0/uJsJeGCSKAcn7ZE1dWADF7zkgYmc1JGdFDrhGVj6KFd7C152to4NgLFrq3mhUZ8+fvypNuqvvehsQeyoYw5MNt1u9DVV80pgGnWBRS74toASQQrqPgBR0bFm4IVrh1wTkY9CUNfAC1Zzs61yFJTqRdrIomXNRZ8PTrzx8N50qMv6Sit8WBF5KRqQ4FXsWm0Ia81vHdZV7YjZJ2TIPYgVQXydMvYEzjZ2tKPsie0IcIFDkIRgWQV+qh94VhXFZtQ5uA95ztkcGKBkc79rVS85a17R1yf6HCwTOkGMJNOQTQKfPP19Do0lVQAlc6vaqw0OfYJmP997HukjT3sFfWqupp08cxfagaWMXJGtmZvmOfWwaM5rjpupaDikNsuq2TX/XQj95LdoSjbasbz7FRjGVCdnZ55P6M4rwJkrBMEIBDL+tPm1USHwmm5vp8gITY9/42NeomlejSeBKt+bmfRdyvhsa76Zhq7XBLMC1tOjnCM6koc/5Rzgp9zLjRy00632eTLox6wjfRjmG2fnF9/Qq8SHCo4Bg8AAG4GGkYYFYoGxgiyWGPmwwLDAsMCwwLDAsMCwQFlAD8/l8OF06Zf8q8vLyyd66H6q52ntcqSHeTl3cjT0TO+Dlno4bytYeLDn4Z0VETiaLuuRHbezyhX0KPrytaEgRxvHRS6Hf+D2w74cB9pEQaDlZMgtEq8uaFZOgR0MXuXC0ahVQ2A1JwdnVP/83/CsxMrqMTXPNJALJ6g5gF59BJ0WhGorybAPOAlOsboGnVkBdsD+RnrNR6+0TJcPHk77cszY8Br38PjwaFrJgt6E/PpiWmclk3WTfKxkEF1okdDFK9+aXleS5+LkxDYC7kD9lxeS7T62Ea70JIHjnOiDEn3YAiet7F+PwIxb+uHFKh6PQcNn1RJFf31PFApWNqaIOUXXbRIXupsJOO9phAettNNWnoUvTjkUssotQQTPJ2NoHjXHD7nWehXP86HjFxk87iwJaTYgmGpdWB2DDvxr8pZ/WPY1m3aiHzrk6FP7czF3CjbjssC92unf0ipA7zXVVswUX+Z40basokkQ2HZDRngSoBKz2ZYYn8T8RfZWZcUkryGeqX0tHjjH3tjNUVpW8QjQuEjeEkGtFkTh+jUxXUe+Vgl2kWQobOXVYKpCouza6FiGsosDZr5Wmk7X9SVKZNVtwci2H6sgtdJytT7XFyLf1OuM6rrUvPXXXRWcQHQx4nrM6k3mL/oSAGM1Vzn/upbVpliDWNfKHeazRTI7zXDZgrnjlaKywpb2tRNzH6yw0WwSM42xDsaHXvDhhZ4EHylzdUDHSddkxis57dgN+/gS7s1DY5eghz49rttEn1WfRmXcMzbgq7Hgi5ZXILXrj/sT9z/SPE8kC3PHMjde8ICOc8GmjlrSSHUPkelwQh+Z1mNBZ8mIjmyKL2Dxv2n3vyxAqvAUcjT92nhwKwAfHZL3Za5pEmqYjwOl0IcOXzdlzNCx4bfriH7LyThLLlaJIZltp3FaXWmvR61M5O8MduL639O9lwAofHw/MO3iy1xSh/SGTniW7eFD8Mzym4fasaf4MB+Rpb66jCyao/Dz9Vxlw4o2LzpC37phfLUoVOs61wr3fPrgk8T8BBLxSBnv+W+Tr9+yO3NAf4rnAKSuIwJkxvN1cr29v97eekft71ycnR0ISy84uz/kDTtOwwKxwJgYscTIhwWGBYYFhgWGBYYFhgUWC+j5nIdojvWlHrjZg4xVZBeAeKWJ/YhyjHiY96EHfQcweMBXuWBvB3xwPHiAX/oLLkEvI+lkh6GjY8dbNO1odA5F6uDVKpTbr72E3ia/vh4aaQOHsp0xHEecpebA0I6s1NOGPnFKwMUGbNbPPmGhSRuJPY/Ao87m4LWipWgBi6PV863AgfYdUyQBHubp1RIVOMBZ63lHbmIUwEKLYEoSbcBwUOYAn3pkTD395PYORQR6SeCQwt9wrTO4gaG5L1MH5lVt9JHcJ08Tng4CVfPMjyo0Iq/r9noLUBaCyMyjp1EQi0ybssAzspHTT6K8eQQ3dkh/zwOY0Ei5Ah8QXXiBQ+AsQQhgQ9e2l0OtGTI9P7nQceqVZESNJJXZhbaYzfzmSBAQBMM8bupX1a9MGrP6rGsbY/NregNywzwCVzTAq9ctCWj3K8qq37iCpw8SKwXEXtc+fEYnwKDABXOb/fiYd8xX2HI9FF/mOkGsqpdepSNw9DmwUU3WFdkr5RrSyiW9Smn6wAuRQ28pGx6afWLPKAJeoWM5BABc2jIWyXv8lIENfNp6GukvnWqc3M98bamHp7yESwoAGtW+yBueaUf+lHu6fZn+HJvw0OttELjIHzrABA77+ZXUTr7A9XgZKa4B/spAm9WxwBDgoh6a4GNv2kjA9Llmovp29PXf1fTi9Mz3O4KSewok80o6dMCFBnOOMkfoaCq6bqLtVH3LdRlY8sixmfd9SFh2acEw1Qt+ebWVOvOedAu36ef+JmffH/jk6EV/ksqKvZYt9QXlQ9n4He3x987WzpYCZCTfw29P/uoY52EB/0AwzDDe5/7tAAAgAElEQVQsMCwwLDAsMCwwLDAsMCwgC7Qn5vlRuz1yX+pB//He3sHjNcs+lFgBJZ9Dz+XaYccP8DggOCIEcnB3KljlQjtpaxRtjL3jIFYCAzzE47zqId5QoinnSqvDtKLGX2Fr3oNcWvfrp/FyBHZKMnhXsosl/rWCDIfJv8y3lTH+NZ9f6tsv7zOakEv+WlkVRwMXzf9Fxo5GCz5gGGAISJCHPzkHex4BTxknka/zyT/BVl6Fga7lNJXDtu/gwJb3yMnqLvChHbgqo3/x4NUgnLyr1YVXvBAUBEe+pUDw/JXPATECd+XkhmYB6Cz5CHqBS6KOfSw//lPTnXZwWS0irUpv2bIAyBstl9rJdIGQrQxScHNdS3Vgi7gkVhAVmPjrn2WrDpVFp8lobxLAJhs2srwCsvyCo47D69UW5QiqDzkkPe0OQpTeduTho4SOM1/VTUc4oU/eAsPKm+CCi33IkScp8oRm6NCfPtqSrAuBJ7Ux98m9t5ZorjS4Hj9dPzvalH8tx/+HH32ove5OtQrnYNo52NdqqQOtJlTgiUtJ+bQreeUO1yoq7ERHBWnL2KWjOiJCySUZalwYLezW+jU3MCPg2FZCVbANGBoJhEEJmyEv1zQH8E2v11+7r+sA1KLJ9aB1QBolrvkaQ/ae2nOQk2sEggp0VMHXlG3nFXeIZmGslW2pOnvR+et/xpFsol7jQhnxan5hidpLUfMFIalDr0sJHqadXmhxMB7IRurHOLC+ZkSPvoy3IM0jKzxX7Xor+ZADYox9ZKn5TWB3oaG+9hnYGhrRbIG1Hd07i/8yD6kXfQ2Hr0tWhMEIy5Q8XqknOGDDx3iSXdoWdeEGb/l4QdFRly3B/QNeO6JTL/kV/dAsmwkHujpyPdF+rflEULje3AcEWciBI3Da5i6zrNmnVgoiQ43tiVbXclzqngj8/ePD6fjooNmkaCEfNJk7yIANS2/pr3/8DTFFxlewwir6yEIgWzp65KU08kFPTaYDXeBpywiUPjUH0NMgpggSUKwAYwZK/zYetWKP8Sp7ygKCQ07oV5ptqSrz2Pvt6d4gfhLDKaDamf/67afPn3xF1yFf9GiJm3jZLS0jHxbAApm7wxrDAsMCwwLDAsMCwwLDAsMCZQGexv3krMdsWs71FayP9ND/sY4LnAkCNHLagPOTO8/tfvhXDRwcBByUvIJoZ0tt1EnA0taXwaMtq3wo01bOSDlv9ehWTmMchMCFnom2U2Qh74/A9vmr+mnrU+qRsccxnAyB3ugPJnAckZXVFfQfHOx55YzACrbpbjh5W6GPfLQ5CCZ6+/oK2f7+oWmEN3x3dvTemlL0iZxu1AkatJFzhC5lUuCD70adAof3F5jkgUmedvJX0QHOdulsGrjgUu+PtEfOvg962Im2wNEW/tLyc3LQlwNZAr9JP+3kwG3yoJ70RWX6Y+seFvjgeCNyaDkoUs4wfQRWYyv0SIpufK7g8ZOnCjSxCf2+Aib1uq/hsG/k01wCx7rijJtXm9OUCYY18szYlCPfLTpEAUgEX4WnSEHFY2km+Na6vcqM/hm+5h4ryV5/+JpBbW8C4W0uQrbkLHv31wWycxD4iv69nMhKO/ckNkWnztcoEwiDtoRxsJGATHCrvfjNZYIb2AEbviIloJrA2SZc7NbrBRngAhuYnnz6vqjN49c6o29gizYrriqw0/MKDDjB2+QF7cjEvYm0CRM6yenflCn0A+OVf5oTodWmR7pr7JudLZ+CY15BpqkD7eAFwXOGSptX9EcOcgJE7MnIV1Chx73Sq8fEGL2A2Vdgmdhrvi5pfKnc07EszV4E7OhLoszfOmBI5PmbRnl9w1d76weLfg7QN8uvGcY1nesamtfCS3K9uy7SHp7UKfdy9X8v1IfAiv8pjC066jtQ9vbP//wvvPPP/Oy/cChrqNv3Pk6LcqqMNCyABTw7himGBYYFhgWGBYYFhgWGBe6yBfxELQPw2N85MnpNY83T9OrRo08eHeztfqK9Ti5xPHE49S6STirp6TtOC44NzgjOKmX6HNzBeeiCY3m4N6VbD/s8mtXjGTD1rL84S155ofYZX7glA05DBYDcYBo4frSVQ4EsHDgXfo+KaJUSdZfMr9pKxXJiNh0ieMeBMy74TQ4caHhgo6urS71WphVk2o+MoAIbm/ObvffEsX0khvbkQl8v7sEZK/amzyo9LMw+N3SAC18HAjobUyexCiFyo3cdvWNWjmAvvxF1gk+NZrWkvGnnHg6dibl43yxodHag3YfsQQoddDFtCUp/7Bbc1I2kU+rgU15yyssroYFPjh0IdNi2bWx6HvNcYMWKYjtJ4Ude41j7DaV/Hq+mK45p5lToBw8c5I3uqdMvq1GdHffAOO4kyf31O115zD0SzjSrSdwvw13pePT8hQiwhxkARc900VdRAL1OZVyv3pKchtH8cU6QoY0NcmMv5Ko90FShDdlV1GdSvbcdQSEHv9RkeakLTlIJGQLC8ZWk+c9dg2Q6ylhdpkn+9hsPBVf44JK4HmI7y9JsBg+CGRwEvFBHV4psxvWn1+S0moc9n+peA6UKxNUCIK3KAVd2Yh6wImeeL7qQrBv0hcXBChyS5yTWlmyaGtbGUvpe0fSV3r71SR+/WgostpP+4CVYAT14Y0P4WTdxg6so0a02apJA+LUaThqKsfkLhjwH8LY7eJoI0M39zTHLFixGllqZVfc78GrOCV8yyywlk0Xw5AGkZBRd37dpYK4oWW7JUbWqQ9/BxqaXYVROoLdkaDZlbjA2HNAUnPfnk00tC3VNGPh63qpOucatxhk5YsPYA/2N4z79GCO92X9Mt02/Wqm/V54bkhR0rx5l7jhwp5z9xUKLfqGbXuYGtJnbpUuNA6+qByerAB1UlH3mpLk0w4go8yF1YCgzdzmwS59kVrczh7GR5zLBc0yZOYq9mLTt71foAw896aj1hXwAQ9KudcfVclfp9ObP/KF/+q3/7r//nw7+/L/z7wquxkaFkYYFPmcBZuZIwwLDAsMCwwLDAsMCwwLDAosF8rTPcxLe2/TgwYOnq/XlIz1ov9xTQMYOlxwfPZwbNg4AD/I4rDz20wbcLYejdyQaDHCk5K60E7gk82ttKYcuzSmHBvlcFgn6cXhCD5y537ALjx53ccA2HQo0XHSDXp+iNzlHeFkOOWf72oesHPtaHQMuvOyUSR7MiuNzriAbjjp40AgMuKyQwDmzgyb82AW4lKELbq83bZswkQ/6PWxwaU/q+2mLzJu6QhNY+jdtAF549nlo0U8CL/yS0w5O8NJOPeXgkrvNzii1hS/tHMEjh39okPf86ecIjZRDo++PLULLSI13z4OAArBJoZV6ctpjG63fnK6kzyePn0u5tsm+X08THcHZcVb0gGuRgC3BlGuCtEr+iAMwpNir0yvt7s4rlPRHRrU5MMOG/3jz+jpmgmMCUrBRbUq2jfC2FXGa7aR+VpA5kCZnPjqhP/M58zg2I6+ygjbNoQeGMsEN7MG0XAIlFRiij0AIATH3z3nTW/KFh4XViaAJbcgCXee5CzYgviiLLqw+ik50varMtTsnBTYy5sBCG14OesxASyEBnZ7u0lvXG/XN/gr39ZDLtUlrAim3IW7XkAm6sc9mvsmzr7tM4Gcet6LVw/TcetrYh+AY44udSbRt4mK7ShU0oh86tPNDzLMXZ9KT1YLa31FzChqQ5iMg+/p4CteD5Wtja35qI0Fr87Bcrc9A7dTLnnL6sTPyQCvyppz28AGHssN2TTbqaXdBJ8vc+quNObqMKXJGjvBQXaT0s4yuWbXdPz+/fF2vNh//3J/4+ZlsCiMfFugtUD+59S2jPCwwLDAsMCwwLDAsMCxwxyyw4Qtaez1g41rKk9uenj59irPxdLW6fOq9wQQht2JL+8Zs8eU4fr2PM6Efrf3L97Y2x2bLsit93e5gvedVGjzE88s7Lkk5BvXwXyse1CZXFTrNR7ATwN5m7EmGH2McRDIATkiV4xyyB1oSvGBUq7r06gtl4ZJwqklyn3TWr/yi571iqhskBLNTaTqGXk7wz0Er5Ky/cGiPk4Rzgg3YjJ/+La342ZIgbEy+p82jeR2IPW+wqalIH+DisMO7dIVByeON/fUqmZe7rAseHH2prASRMNdyEknb9sJp7+io/cb2VDuSk2EQ5dgg+vb6ya20HNgPswIHz8CQE+SIrJGbOuXQhE/216JtoYEdikdg3a8AkL8Up4BHeNHOHmDkHHFCUyYvnehvAQmcbtmgwiultgcNUOjZXMVDvbeS6akl/KNTcsbaNKQrCZ1ItKU9NNyhU+atAKYdXSfEmhAamoxzzUsAEySQoFZKesvRf35yOX32/KVWlOnaAAw9WEaEmqobVAX4OGETXaPMPzXy37mBKeNtN5hCqPlTLAWAfKwE4r/mrJfdRV+1XcNbuROw9Amef7pBSCwFLXQNvPn6A19aAPNaKDznL4VSNsOFlG14o1EzKLooCCcdKXlFm3LPIbWTsxKJ+VCkC95zVhjYVhDqgwvzsnC5H2UskZvxdGARHVqyBu3acACLIJn6wDNdiLkFW1RwBDpcE17KZomZq7UCLnTJoQd9El+1rES9aFPPPEqZnLTIjdFtcuezXKJnXIlXtpTcGqsWg9IQwY/7qwDMWnZUeZZD5eJRcuW+mfmr0TA/xpgEFPDcaz1pTFatvl7hXfSlGQCWyQXdt30Nwtv3lcZX173HUzJCV1XbkDngRVTAEiTWv9OTl9OTZwoaq8yPB0f7B6bF3wQCZn2ClucUjcjGnMIGSubf7p81l9qcoV/qspcmZtuBZgLcokFCb/qY+0VPDdjQpAsP1bG/x0Vl36PU6Gu+7S2HfS2HCAIncq6Luu3B3GJFNn3AoQxyld3FHxl01iqyG1ZonuuDMVuHh/f1mvLxQ12DLRVUaj9SXnraED8S/AD6J9ECGeV/EmUfMg8LDAsMCwwLDAsMCwwL/P9mAZwInva35dj+X7/x69MnH/7gmTaG/1gMT/nlXf32UXjtxA/p6sAR4KE9B3D8sp8HeRwOkmm3nDL9aaeeI3Tooxzn81V1cNLf41OOR0gZOm4TkVqtIQdJHgixtbRDn7KdFPBbSj95gg/QQ08SThc41GuD/lpNgFyRLbBeNSNY8CmT58DxCn/o0U4qvqUndRwlgnBJ9NM201EHZdr7lLbQoy8wyQOzmacffZJ6O6UfvKS0kXOkLzTCYxMOfNo24dKOriT4k6AT2n0euhkDYHu61Enpjzy0AccR2pt9qQcueU+PclJopU7e00h7dAo9YJg7jOSLl6fT85fnYJZ8WiF2rUAssKQZl0rGQV3Rz/0N1iDYDx2bHSm7TkRE1zershwcwfEnmlcRPV83BQsVsWJKgKsAA6PPdeWPJah+qFfeHj44FKo+hGs6izzg9gldN4NUs24iT/Jrem2802c8qULeH4WxtKcOXmbp5hyz/I1O5hk0SYhQ9Lk2K3gTGZLTn9VgwQOXFU75Qmlg+XKtWmf4jBPw4AIX+YJD32YqmW7r3sOn7GFquoUGuMwLYDh6mQtmaQudHqbKy3Wo0fXfgwoOMS3qftrzW/gs9zjo5MDu4UXel7HtbBONwcm5vhqsa4DVg/usHtOE1V8Mv16LXvymEP3It7VvY/gTOk/qbU9beHK7IwCb+eI+R8TKZowh8kbm4PV5yj1dSWV9N/lGN2CxB/XA8LcHWaCXA52SAk+eObjWKjLtJfqwCxZ6GgRn5MMCscAyk9Iy8mGBYYFhgWGBYYFhgWGBL7sF7P39aEper66m//a/+a+mf/vP/punz58//USvwDyWI63FEFu7coHkaeCG6DFdNL03TnO0ysnhAZ7v1FXgxhz1UJ8EDKmCTZCCyOII4RDgcCTvnYDEZ0yDgJK40F98iy54rsshx7UJPitpWPmG7Ha0BG5HQkp4JYOcFmSCdwmoOr/mV01n1S1qk7XpBH02hi7nBeDiS5CQ6IGwLA+BDuTCufHm41BEd+SRACtv2oxDRLBLzaK7J5mhg961T5HwtTqAACVA3qidgAR6RY8aG/XL5jriTKGjrCF2cgwbLHVLvDE+4ABDP4f3RBOg7d7y6BK6tiE4TcfYPf3hGX4Z/8/Ba2Zty+ENL5zu+IHQ5CgcjZ7mme1r5oJkfDzGeg2VXLZJkmi2dejyWhfHPC4KYqAt/TnATTk5tmGOcdhOgqFMiq1daSfmE7i+bJAf+tIpezKZBnJqXCSCaYQeeOjI6sMPH306vTy7qH7mKEFSEHStslqLIME2QVt4kXDsvd9d6WCa9DHkzAvhZH4YvOFxPYuJ+WB7XyWegJJRPKHu1yqZI6prus3XGHTcJ3hWt+0r0K5vUwhG10BNtbIFgErwYl4zncOT8WWs4MwxJ1bstFU72MzjQZPsk7HxnJ8RFCP3XOA6KRt4fOiXrujBYfvT1pJfLRV9L0DS9cuKq6w468c8PHMvWWkO1hcjY7siSHuC9Za/jTP4pFwHlLlkU6e/riHZAwVk6NJDQM0yoQEuiXoNVWgvsOgZ+bFZjmWuITftZVvbiiHW4HCnhbcP9ZMo085qqCTkpLp5HeWaBdYB38YDe7DCbpFL/Roz8Nn4Hg7olC88wif8kG91dT1dXJxp9RgfQGEfTIJiOjR4ZcuiDV7poLGQ/TOe8I8Nox/1aqsJ668tMxa2bV330OIgoTM2Z+MBSTsf9C16q11wmlVC0Hhqztc4q6o2Dnh6vDXnuDdkfGocak5RJllG+HU/lMSGMx3dC0TvnsDfePniREvIwEVSF5S1xFTxdEHf0jldlYPCMdKX2QKvGvkvs75Dt2GBYYFhgWGBYYFhgWGBH9UCforW07kewq+nxx99cP6bf+/v8iXLj+XoX+Co4ynoQR24lrngh3acHxIP63G8AOWhnbw/gKO9f7CnLTD09Yn2PlEPXdrTn7bgh17gLZt8hMBv5qE143VMQzNNcZoSZPEKsfI2mnPbIOVk7rVgzIFel/Om/bKl8XC1FCiANgcPqnEIE6wj5yCQEHlxpihHplneZqfA9f1IE7i0NwlvZX1feKSNPOUg9W3hS1+Pm3L6wbFDKDjKaSdPuZ9D4RW69AWPPCm4tKWfth7G7QSCCC42e23vau4S7VFCrh6eemRNX/DIOTyvJFPq0GHM+oBA+nCOUw4/8j7BnwN8eH748SfT+eXKG5LbLoiK7FpJ5kAT+mgu+RW/1gcP6wocR5MvuolDz7KCCti1tRrfl13ZSsQsd/na6lC99K79ztjAXqKKjyaq7h8H2nfv6IBiBb2hB7yDSspJ0TP2tW5qj33IA0ceuOTuNAD6FSwrQ7u4zWyD4PQ0Z1tIF5NpeegGljpl5EtbcnFrQY/iH1xyeALXH31/2iMHfbSFT/p7nM1ycIGFH3XKaXdd6jkI1LX3dIB/VYrN0get0E0bec+b+m0YrtVlLloeB4mqzR9gEN2MvfHbGHIvjGyhiR4rjfWF9mvk1UqtkvJXgsEjsOnX6gk0Cdf3WM3Jrfa3CRhB+DzTazbp6/AMX/LIRgCe65fAp15n9A8YgSXvaXD9Bzf4THvakoLjQLE6wefyIbnc/lb5/t/mHjgc1k3wfUofbQI5lq5f/fTTT99RlW2moNyoz5e5mka66xYYe5Dd9Rkw9B8WGBYYFhgWGBa4ixZYnsn/YdrPUKzOkkd1cXpy9kgLCx7pYfzian11dL0SyM7O9Y0cDh7GdwksKMWRj7PDXlvE03h896/h+XVaOL0TsVnma3G06fHfdBVqs7OLY8HKK//6r57tnaLDXmJ4AnGkjEubKIS2CdGidg6SSqKFk04dJ6wckuCzGkkEbuGUA16BHe+jJBAHJC54zae+5HlwoIiAEo7ltr64x9cJvWpA9AmSXe83u7VVUry16hUP3UoKVo2Bf9VWxyAzetKmLWa8cgKHC1lZJadXabx6ag4KEChwEEZZsyersqy/VJ51xKgtpY2clDrGTzl5+qlvsbKl8TAi5lSKnVnEQz90+NfTMFwT4boJ71f+RBedBCw1WGXCKjLpLhtAFxq1L5DGgnLNMgVixLx8XzvQvArH6iXzcQCJeVPzyo06QatPqZPDkxRbpy+Brzi9PQw4HMExAWhohSD4xmHlDNbQGMGedqSgLytR9MKY6TC/uOQ+ffpyumS1lf6pR7iyq1fZaGWkXjNTNKpWJoq3VzPiBotu7MU12JjQMW01e8C3xgo7yeYmXEWXVZRg1a5+JPUqK48PWshOoKKz9OHjAOjPvmUPH77h4bgSLDy43rBd9BW4aVFnXtdX+SoYYRi1o62YwBVJTIc+IVo8AiKef0imdka34pxVV3P1qw8K0ZfVl8Cji3OIK5UtgKsxVIvbwfMh3Ugr7OQk2aUTyWN7zTcqsYXuSbaJrlvx8f1EtGwrYAvFeB4jUYcksJHBndgcxlwOyrCZE3AqML37uRZcT3sR9Nc6hUMQ1eNCm455xSsCwdiBH2WCLXo01xwtzsW2cGU74VlfzeWkwNcrqG3lJDozH+Ch/zAAD7nYB4357vuDu0TXstS1ZxxmgFhAU72eD7anDHFxdTUdKwJ7pGWK8CAwRk7yHHGplRln3QOZN6Q5SK0mbIFssK4+ytgIWjUu7lJbVp+tfb9mPNWvYFzpqICY9oh00r0evUod5lrZi90mbV/Jiq2pi6jt4fsBlyl8Ja+wJS7jLFr6e8xqtt12//LfWya7Erpyn9Ar/luaizYAPFQ+OL+8+pr+Jn9NA/ahiCiS7W4YgCfxmtKqj3R3LeBZcXfVH5oPCwwLDAsMCwwLDAsMC3yhBXhabh6Es/M3H77+Q7X9UA/k53E+9OAtv/L6hjrOIQ/jJOrlKOBclKOQvJydgqGcenITaCd+ne9haA4d8hyvwu3b+jIy9nXKRbPo9fwp09/Dhyf6FV5hoD+a8moPXhZ9BMWWgKFcINXx28CNrTAPAbM9OUrVj88innJk16v6QhuOGyskCJjxlUvkAT8BtJKgO4teiwe5EX6k4EWf1N2pE3DoQYpugaWNcq/3Zh/1HOCnDE4PG1o9j5RxCgMfGwGfcmgu8DW/vPG74DbbU3cQpkAhZ3qmKZlpjnye+J0ewKYPWsjGmJJwRtPnhu4EbGSmOXJTpo8QTnCp9/3IOuNqIOG3o32TCDZ//OiR+uiHphxxgmNU9Iolx5pNuTV/KsikMSUw21L4CVE4y1gRHKq+WuniYJFA3AZtzUX4ILVXAIFOu44t0+94yIFHnx2i4pKPwNXrD17THJfeuaWo3TqZXuHGptiXBA3K5KRZ9tZHG3OVdgIlJPPV/AmOCi4Dw0F7ykZoJ9oc4O7qFIHfPJgfauR8S6ZcN+5ofZEP+ugHLezG0csTHPLIR04Cp0/p79tSBvZVdHsasS/5F9EKHehGDsp9e/r6ftqSep60hS/tHBolEa/7IDTKLsUPWM2u2U7gh08vA4HYS83NC815Vo8xN5lvznU/5QcH7scEKHW1zfMptKBLSp38i46MG/dizXrDEaj3vnIaKr8Cr3tzxjY0mQPBjY6pA9OXCYyR6lpYxidwdf9PwLHGI3YFD1rACB5CvpDAVcBMxrn5McnyY1u720fAtgQcK8FTH/kdt8BYQXbHJ8BQf1hgWGBYYFhgWGBYoCxgp6U9I8t1i1lUwE0hXZ999PjjD/b3dz+4Wl2zQ7gdBOHpmVxrfvSAzZ4x0CG1X7ENo69fqn7odp7ZG0i9fSUnBm482GfFRNFQcMjOM06CAjYEj/RmiNyXGb+e/2f5RLkCDtCL81dMy+lpAgi/ghvInCN95VeonWUeFhRHqFb8FD+d20oJr8gAcXYuSndeKdvXnmE4OdiBg8CXbSyakKVMP84TK97i5Oxq1Qkrz3Z3z+T0XclG+hLmuRxqBcpYMmJ60pPEOCF/bO5GnWiDbmjSTqAxQQQMbhzJgd2Rw3Ywxa4+61WUwTGcRKGs/7d4R44ZrsmGHPDBJS55C89tjSYcNH2IpxQPBtHjXzYFTz00lt4qZwUObe4XD0VqvfLEumppjmUpEoIRf/Hb1viQaI6sbshJvMCnjyOpZC8b0B696KeOPimTR7/kpQOzSDQVnGLPJaeWY6H6V+3mp7GBjw9tdH+qL1g+e/rClmBvL75qCZ0bveLFNeLFnrre1lf70572Y0J878XGKkvpVXYS/djTrJqOakMPQVmsyNsqxnEbuJpf0AA+a0+MK1JbmsNeoCK5kHtLc/etN15n4LxX0h4yKXCBXa632FdPmpuv9GEO6B85YtBOP6mCH8JjqZGSacO/iU8b8DAiQ2+Fz5h1Cpo4VgBIg1FB19M2MJp04GWlYvQysE5Z9cZ8K/q8VofuEBMZlZFRcRofhCa4NplmXIfcbpBVhuK/7WC9hOcVb40GbdAiiFj3wtJb4RIzmu1kIqLJfAZe3R4XQfXJgUzLolblW9y3+MFB/0jGbfdCaGuWuSf9BtIpcoVH2WBptzgiyR3bMI0mLTVGNdbYBdieHvDee0ydfmVREtTqwoZrwVUWnkBb4npgxRm2mqaL8yvfr/ly5b6CsvBgvOGTA8SSRbmwci8qgqLDYDb6WIjUpl3xXZirXXpqaJDbe0YSFONvhND20EM59xrdvWea0COQRsPefE238RVvVqGhpO87KiMOK9SMN/9IJGzGiU6lCgLKFqzcribJpFHg2qRFcMsq2ZtDXZVf393b+vrNaqVgmQEkJ5OiFMYqGWMIjHQ3LbDcKe+m/kPrYYFhgWGBYYFhgWGBYQFb4BUPxjydc+h53O7q5S/8wi98IOfhB6qf4GxwCO+GB/L2UO4H7PThdJRTIgegHtpna8PPTglMVAYuiToHyXBydsh5+E+O8wB+4GbY1kY7xyYMcLRBK4l6wVXO65C9PKERXn2ePuSJc0I/QSeCYgS09vQqZU+P4AjOI18HxKPmF38SsPsKeLDB9NExQbJFDmAuzi4Nmy9k0kY5iWBAgnbIZe01/uMAACAASURBVFe4OU7A9DojI0fkD420p/5FOXBflDb7MvZpT24Zu3Ho23FjSbTlAJ5EnsMN7ZS51sOBG9isMPNm6cIJP9DBDZ/NvJF3FnppAy9jC5/QyVylHnkCl5z2yECedmgbX/2eU9hAqjMvn7840Rf7zuagZtlW8wibYDJWkylYdqM9mVaaGzjtONViVCKTC1bMBC8EymkThOWpKKV5GEn0RN2BBUeA2BBcZOKoZ16Bm5Voi158POF6un9sn1zBYOnZRGGGMqK8KubAADpwqD0JOm5rfbT3No1taXdgRNhZheOADPq1ZPkaPZro5xoJfdr6cuDTTk7iGuv5Akdwra3c8ZjRj10wvVd8IoaHYblPmBjNAoJGEvLfrtc1EL173uBswtKfNvIePu209e0pp5+8P+CziTP3oxs/YGgcQyewmRvG99RjHhHyIyjfxkYxmrLVMu7AR5b6GurtcfIr1kLnWj474/carcBlL0ePJ0EozW/4EXQSQ+6psrzl668z+IAbXQh4pZwcCOSD54qxauOo0KfH1uNX783OMgeX+eUgWnuPlj+lmSfMC+PKDrEbvMCt9hqDtPk6brLQXza+bRdgGy1+tNrm/lD8pgN95fOrf/SP/7Gv/rGf/Vn/WjVfhgyeEnxHGhbg+hxpWGBYYFhgWGBYYFhgWGBYQBbgYZ6jPWDnaXlbjgyffZx++MGHT/b3Dj9RUOYFBtvRipYtrQQBHueIr5zh83gfLD1s02anTrB2pr2CAWeE53HcZkI6lW4FUXAum9MAbfx1r34QBs5O7VkjPuDXs73pQYmHfHDiQFDPQRvJuWRJO7nbkJ/gguiyIoBEHys1atUYj47Ck9MFb2TBamJonsCySAD+6B39y7GVPRwOqP7wxOI4MJGNlWfHh0deRXZ8fCw6RZv+9fXVdKU9puToyCk8cw4uMlUMs3RCKm9OLRvizBE4Ycsd5IHvZprbGBfsjl54l13yOGC+blw82DOMZk6jbViVqXPgEiNHeaxV59VR0/I8ICTSDkQAR/yhQyKrInXmg8YEmoIr2xYcsOapKqowl3nfqgIO0ksTiVnHK1cOpmiMilebL7jXcnTDVwPt+kxX/BiH4MCbFPjo7UadgGNeZ2wtm9q4TuKIBxbc0MY0HOi6Lfl3/NVVVonsTh999InGni9YMsaMe9NdDTfa84sJ6KEDgMmo3HOXmJad+BbEMAEMJTujh+Hl8hO8pSw75ag99nRtBBbRNKCsbrzx1/PAl6xGg16NHWPAnDs82J1+/Btf4xsCosHqFl3H0m1J1BlTxgh7SkZfn4wFZc9wdbB6rLD6fQbhy7XFHlCxNRjME6uiPvIt9XOdeMWS7CbpvR8Yq8E4IM1qsZSpU0ZvEuZrcZDF7rSLLnNsHgt4q07i+ry80KGPKtRcKFr0QRd5M/b1qh6Cip5oeB83aGMr5ixtbf6B7/unlqlFvuW+KhrtvuExgyRsZagSC/nCe9EPikwFRoODhGyszK37r/rEP8nzqd1HCRxdEfAR9GwH5kFb3cY8MC3kaDjIgE3IOUimzwoqZBY1rlnGMgf0uf8yWsHj9cqyY40n10WuDWC4l68J8mJX1Zfrr8aAa3G+/0i9eoW9YKFbASYJJP1YFYgJVrpA12utXEO+dph++3tE2bCC83yTTtCyvhpLchLyVLnsTZ2x871L/eCw1ycsgOOolWPqZIxbIFCE9F/Wafyhzd9cXaNakLelLd62doX55re/9ZNv/cqv/C8H/96//x+IuedoTVTbGKyR7roFaibedSsM/YcFhgWGBYYFhgWGBYYFOgv4IX2p8wC9tavX/n7j1//m9PyzTx+t1pePEhyQ4+N+HtxpA5cj/XYU/KBeBDdoz/D00mcno+V9G+0kHAbgklOuIJG7jU8pdHp+RaNktPdSKKYXHPIeJ+XNPPoltwPXHB9kSzCKlQvARH6ceVIFAsqhv5QTDX1sKM2m3T2tINPrcXvatKn21Vn0xhlk1Rg5elOOriaM09RslTyyu787xYZd0+dwQwNYUuqUoZsjffQHljaS+dtDX+rYhHbg3V9dPm+2bcK9Soa+LYEPj0mji0yBIdRACt2UyQNDOQm4yJjxBq7H79vB6/t6fPDCgzx44FAOXeYPB05wBdNwmremx589cUAL2Nsy4XDrumO1pYJWHGtFpK6vdL0QNIMvTJSC5xUpTQ/aK8hKqeYnQQVFFxyMoM3BMHnqoZM5TJ+Qb407/LA5gStejL53pP3INF+xvfkTPUiCB3NBeZ+gkQQt26oFAFjNQ1vp0tnCTv/tsYFGYMkJcsUG1JMCQ1/66evrPcwtvEVUmaJ+HEhAg/xKQbIVAaTGL/aB9m2aJXv4xwaBS528L0eWtJODk/nldpl36efHC/bPuz0HN/WNHLQzduC73N3TGAsSsOFb+WIU93XjS39ki02gkXZy5o7rykk9HyJv9BFs4wcDEnXut1w30NalIBqSSeLBvz9ic15tpJ0692GvEFOdMaMtsmWW9G09DLz7I7y438M/9xzkdB9/KxTQwv4FWwE/6wRQS9QjH7wpk2hHR8PrWqoyoY267gTrbQ/UgOgSlet2+3W1v6lA5tGf/MV/Sc230ybv272jdlcsMAJkd2Wkh57DAsMCwwLDAsMCwwKdBXgE6o/qwg3xUf6IanEL5Ntenk//9X/xn09//s/9Wy9evHj2sR7nn/KwrgfvXeVaZWZHw0/veZDntUO+tuVlBHJsE8jCWeAo56AcgJKgHFmzh548WdykRnt2DsBjZQnt8AIGrzf1V8FHX/qSKJdTULbwXk1asZNEP44HARdWqlEmyU2xc1N7mbGWacGBHgdkcNRST27biKJhRM+y4kAr0IUTY5kk4r2j4+m1e0cOksF3T6v1wAXm/PRsOn15olcuzx38iL296kq40I6adpwkoXyxot3kQw/3IWuTgzYSezwBn/bFTjU+BaV+xUbh5UCO51PxoJ/2JPmCTmmjh9VH1JGdBI+UaYrj6E6NMKsw1OqjvnRXYxecgrvNN22MWBs6NzF+c2qGimxuZ4VLm0/IhRPOAQwH+sKXsvsbsdAIHH0c2JEUWYPDyhbNJNMpElqtIrrAsZrIC8CY5yzDISCg7LnGvQIbRRs8v/Kn13FR0rThK2QHtFhypdcu6yuXXCsyLgY2oshaP3RkzBUQw9mWVN4bi2ATsLI9+515BZLgomf0EICoNZoq0c7BNc5Ya53pdCDhCXiwNonABfCsvqkVZTVuCVxllRnz2XR17bFSZrZ5m1pcf5Di1VmkloC2dY2LqkolCwhwrnFHt5pDBvHJ1x5jroP7llfBSmXqjL3nw0Z5boNPgpCSpca77MHqsXULZLMyiUFkvBR+0S2LlWvYABGW+xf3G47YWdThIBByNJVMGo/Ss2y9jAWUNFEkM/MEvUnpNwlkgIpyaMSutqWEMV/JWJw014H2HK650d8XinbZN3xC1+NvOZoM0ER0Hfn4SnREhhor3Qesa9nPOjqYWtcbPFhZR0I/grrg8XolcrGy0Ht8SVFE5j7MvcSruLC/57R0VJFxJsEbbmZDEFOHP46ieb9qB8G5K9mccdGCLB/Y1mNqKpywqWTjOmQecH+UDPyERDMJWSmv9DENjwmr7DwowAgeEQXDgR0IooEwz0f6oCVb7upg30/D5po2l+UkmygOXp3KxG37wc3q5vjZMy8CN2CNQdl/wRylu2qBulrvqvZD72GBYYFhgWGBYYFhgWGBzgK4s/zTM/hm0lO5ntP15PTh+++d/Nbf+82P9FD9kZzKSz2A8zzlZyqcTA4Sz+R+4G9OmLBdT5+dA0PiT5RjUa9yVWP6k0MrATUg6qG+cvwF4AJLf/MJ5rb0FwzOwBKgSR94myl60B7deN2IoFjpV54PNOjngwTibueMr06im1wU59DK6gZWiYUmgcPIS06d12MIkj187Z5et9TeOi3YBo/SXXC8bnl1PgdskKHsVHnKZtROwESn6E2eFBrUo2/GJ3CbOfRoiw7gbtZpwy4cOHsea+GEFr2Rt/Sj5fMJHsgTPMpJaQudtIde+t0u57JPfV+vBzDpI+egH5ocsU3y0OzlAh482kKDPDTIgQlf6jjAgYWmKEwKX02PHn+m5Zzy+tVPjnM9w4EjOnO8Fnk1Xwje+PrF+aYf+gQcm1yRmRxYy4F8OojSza9dggNN2qHBf/KWXKZftwDKu7v75rMjPg/vHXtFW4sFmEZs1tsKPAIrfYp+5LElQQJgHbJRO+XqR0TJp0ROexL1OqqlhwsMOfeZdktr5aUXeqEZeq9qA8P7Dypws9YrclzTJycnCoRrPJoc4EX3jD19s44dXElQ867krrkU/E0ZgC+4wnS/xo887QSI0HVu030teheWhp+Jo8T88yb6+iMQ+cKTPCl9ZcMao/Ajz4HcBStMBZyKFrzqHhF6gafely2n5OWHhUu+3qoETQJGBMmc87eMaJzTcu0RdOKAv+/Zyhkf6JOiQ3La+3LkQGZ4bh69PUov2Vg0uIfvVHTY5eAZRnoHr3DqByACncgY/hZQp/w9IAAIfGQijh06wDad9LZx2UH1BwcHhw8ePnxoUoJVE5HDkYYFygLjK5ZjJgwLDAsMCwwLDAsMC9xBC+CEfHHCQZUr01yjyni89sP29s2l/ImP1pfrj/WrPZ+N37+R46WHfS0K8muWApUjtkHeqzbkTNBBcIQH/qQ4U27yEz+OmpwS6OB8Nccq8OSFX1yQFLhaOUGvHBc7cgo0iRdyl9NQPFdymqodPSWLVvK4LkeNXDu2QESp5QTTqLHyojkaUCqaEk+d1y2wUDbQ18z0eiS/8PPKj+HoF1xZtQImDkawRw1Br+aiICsHjh+8eMXy7bfemp48eTKdvDwTjS29rnUpG8rpvpRzqCAZ8HzJzK/UlRHNc8XKIetefFlvgyzoiP2ipk0sfdKuohOwBLP0qQDjRV867bC1IA4rg7AV/cyFmM2rG1RvJrMsllVjbFsgGw6j8j4RvCxZbrcX4YUXWpmn8K2n6LK/kNfNSBbbFNrEkzbm3MwP5e2gK2N8kAkW0M7caQqxh5Vlld6kol+BEMYdWWwjObXYwWqpjT2TCHiW7szt4uNCO5XtJKdIV4i5OhjOLe1Btq2PN+ijptOjJ09nOsgJTXn7DIgAhYM9VaboFWQ7zNT6wl7FHlSXXiQ2/WfuCcEOvOWFDoCqcP1hDK/oopPVLBlP1bfk8KtVbXBTNwIRvGOu6/VMVgkdCGZfqx8f3L8vdPES3lpBIuxB8MV6Cw17gU7dqsCa8VTgAjsTEChmyQBGViXhyNrWWa0O0KnRXbxCxxpQJ604WrO3oIUmq3tDdXJuwWfLIjlggamgj/5K8EEHp2IhTrzSJ31sS+4nNfa08UVark2u57PzS/W9mB4o6E1gE3T0Mh+CnRoX3z80z7ifXLV5i0GYv/BBjsKUGBp320/iwJOvs9p+TT5sTN1S09/GHfmbBtZNdwSrw35rjLHhKKrV9MgNUSfaNYriV/cFAlLcD8xKkOjtFYi+Xwpa8x+5CRSWPGaraVL3OWiLgmzBfQk50VOzr42D43bQbXIyu20H6XN+cV4/KGhs93XP3efDJur3xv4evGY72Zv95ZhzsUNWEWJrErPE8kkg6HNfI2c+SlnRlR7KSbSXvtfTnuQFzyvFpK6DYc3Wha97KCs8lbQVmHO6K/hYY8Q+g57j6vW9Vfqv9Hq079MSADp1n1IAUHMGfrElfbQxd/hb5pVx6kdP9emyXGBVPtKrpK/v7OwdidWZumUgGQf6+n871byQRLebR+1LbYGM+pdayaHcsMCwwLDAsMCwwLDAsMDv1QJ6pA4Kj831hKxN4rXT9umbb775nh7I39XD+xkP3zzEy5FlI2Cex8sB8QM6r8DMdEyPfo4k+nPgkPNQT94HVYA1DJEOgg8bNBZqRTU8yXte8nIEsK3AVT0Chk4cpsKuc/qoRb7qKVPs8t2CTg7KzQ7Wwa/8SFwB3cLfxKFOAjeJcg6CTMj34MEDO9txtOgnOMZrljha1EOr5wFNXkPKq0jUgSVFr+Cl3Z060R5bpi15bNb3mw7RjJYYQwfAVAe+gosa3zYlwA3v5MFFltAOL2CKTs0h6oELbHLoABsePf2UyXH0gSFgkVT1kq2n1+OFfuQJDu2BCz3qyLnZnn760g+M56cDBTVPr7WfGOP+Qpvzf/b8uQNHPZ96fVLyowdzu10j1OUtmw0b+EOHhANPXy+Py7RzKJAhgQpX9djfyJwIKEB7M5lfm1uSwwE4WfhIQaKDwz3rCArOPPxicsq53pEt40ZwLCmyBq7a615Aee6HbtMNm5KYbwTroEeMjuNKgWnqOYB1gEE5K6XmIAyytQNaryr3bcCQIg+yoO/e3oHlOj09n16+PBVfyaZxgm/khT9lUtro7w8C1tCmLQnYz42ROgMXWZIDDxcH0JRDa+mr14epc4RP1Zkzi3yzrASAudcpRe700QZubBteqQNHm0gYrvDLJguNZa5K0qIn9Rmj+mAFX62swBi09JvEbI/QQIZcq8D0BzJupuhODg3kIznw1tqoHyhwDV2uT8Z5p+2BBk5405+D+wzbdtLHB1nASSCz5+l5Kh3rYwDFvGiUbtlrzbJxzStFVld0avNpS7py+BrTK6FHwnn7/Pz8rbpZOC6YyVSDGwIjv5MWGCvI7uSwD6WHBYYFhgWGBYYFhgWwQJ6G27P/FxlF/qUcFFZrbO/rta69k7/9t/7v7/7MH/6j39UD+6kdHa1kUJmHbEhqzYoyE23OalvZkAd4Xm/BMfBDuwDjKO/oQR8nft4sXGRwAOQSGdarLnA8xARaOAxFU7RwWoDsnBcc0PrVvRws+MwOtuDkMxR9lUn28eT8i3K1y0uBv/wL96OU5RG4ZRExutADWehDr/3dAzXW6isc2j0x3tLKgx0FKyw3K3dkE8reCJ1VCTqoJ4HHHjvlSPIFtpvptQf3tKcbX7HUyho50zj3L1++NIw3sDaZcrq1KZyCAo2edJo1UFvpgFV/f0lW8T94WObyz0yMOvRxX3GmqXNgowLwKFVZ5wV+brItPTeERwKGFLkpY++k9BPWwNl0j1CutYKuZAkN5otwhei5gN1jGLXltVtgernmlWSijSTggsY+UqZPoxKvc2mU57FFklqlUnOVgBEECMqhH7i2i+YpZVbeePZJN1avENuinbHfV4Dp5LNn07UiETvsvWTb1hyCt1dzaU74lTI57cx96wgRjvZqlxgSocI4ENehXN23Erb1eFXHPHbAQpR+jCT8+ZVNj5H6m02whMIQJlsre0CpucG1QBm6fHlS/13munMIT/cH9OZaAk6amA7BVsaXthw1moiido+sQIVPCj4rl1iZlBVD/touYJFHuLqITIM5vbV95Vf02kyRfMKFOvcTyaJRFQv0p04TLaTiS8n3A8EbT/ZibrGajPT82UsHt+9rVd3h4f6sC3NH7MtuDA1yKXE/XLXgZt1nBKMuzxHJ0cCKjmxacwZ7VKp5KBxENkmYSJ+NoBad2CR6s7CItATFXG33UF1tzAf3S0vwBM+9kvH0HaKNA22e+4oy1VyqvHgVTc6K4rTrWgREbo2s2BwxRJ892yyL2lhxhZyszPO+Y16pW3bnB4M96wkd4UivzDkhWT7k4McH8tjZQTDzKTrqcsrfHc0+w87TXzYMPmKy5xgJui041fRhLpZtfWVLHtseJCeNO3ZTmXmKPNf62+NXoz1oDUwCbokOK5NzTfieo3b4kTynG13PA1l+fb3aJoBHn1bAHUjjd8TrqwJ/LJhzrmHlWNcWNyGflvm8tI3Sl90CI0D2ZR/hod+wwLDAsMCwwLDAsMDv2QI8WC/Oi1/e0QP09o4fsLXJ1i//8i9/T87e715cnD9SEOYP4LQVfOERuOkDGLyaiCPBgz1wfGmPenjgTFGenQ2Vbyf6y5EBDvkWnuUUAE87KXRckbMgyi7WK5JyA+Y6jghOmbsLXPR51Sd8WiPE5/5dAhAt4VThrOCUVTBLvKRnVk7dtmWwSlbgvQkzq1rKSbEzB/6NXlG7uiqbBItVaffu3ZvOTi+IztgRY0XKLKtk9Os1QkCeeQwEW7YpOwBP6mWjPMtgG7QAJrBNdyO1EzRCJ3lPT0hzuCArJPC/sD4JnAQwer69HI3VzIc6/Umv5pveBRY7yLwLrnhbVqSRTOU8s8qj5qGkuzW/NuWDg3k3WSKTA1wwsskkZ6k6jwPjjc6k6EkZWpnPu/Kc+ZqeZruAtLpENMDRdnbTx4/1mq1er13vK1AqPsEjWuJXJT2RCSg0xhAnUddBIIFAqh3viIcDzoowZaWHbLBVzrYajEecJLZmbnqFmcnKjlz76EyCDzKIJvC7kvv6cjXdP76vlTYKAqzPfW3wAQL6sSspOW246Z9LXE+2dYXcCA+QCA7s7EoeyrwGrSJwUOCegr2h6f2mEE3t7FdF8JlE33yNqJ756BV2GiZEKb4l01pBC8+ldi8yEZ2QH1okj2PoY1ul0ovXrcv1ZIzPzs7U81L0X5u29MVa82m6c41kPkQ+8xVd7q0EipC1NG8623ZpWXiGv/NOlmWu0/OPTmWHguN+h078s72b7qESWzAQ1l0BXcM3GROo9P2vjRF0Qmvmxb27o41ZPQ00H5jH1wqO8TVfXqsUJ9uE+UAwihHe1bW9LTvx447tmPFQjqmv2ziGb+QnL771d0aQxkdvw3KJSW7K0Cdo5SBc04EZyGWQH3rC3/OJIJeVgEfmV/hVjl3QtQK5GNES6dJDt1qxZt6+3lufytii7JzrhT4u0bpeWn4gmK/rb6GOre8q0HtefxfXIp9ryQyNPE53zwIjQHb3xnxoPCwwLDAsMCwwLDAs8AUWsMODYynHYTPpoVr+AZ74av3+e++dvvONH39fD/IfCO6flbeh5WM3/Cg+e2g8bOPI4VDj1OHQCaYg5BnUg3w5C+FHMIB2Uj3MlyMGLR7ieX6nn3pyyms7x+IHedVDBxycG6+qoYQ8SqzUIIAEPfjstPZyWPrgnexgpwqPSHhy9HCG8TfMt+1tjOLXWu4QmehnDzIHX8SPFQVFx+x1KocLWiv2YxICpMAvCRWz0BjwNTUHDySnHWJ1Prh/b9LrMdOjRye26835lXNpYrpFQ7o1VtSJaSTASHPk7MvGwwAtpW49sZXa4xDz0QH6MSD9FE1TjFjdRKKO9au98hIK4LK7dQsMg9HKLnQneJBMa+ZZ86BWQMVxlb08d8uxZT2EcW5NZ8muduZiHP1apYKtJZiFbDoJCt6Gow9DIkdlnmdi0AJs9CNTGwk8XNGCf+yzo4mCzkwHxnzWC5oFVP0istaKIey9rf27+EjD3uE0/f1/8L3p7FJzRvFZ5Iew9UMoEnJ5sFUg8KBrrl8httYr0l5pJl1w3ucVKuBKrtprrKcjHiIV2QCDJ6xR1F+2pCgLWQ4UK7EQUNdbrRR95+039Qqc4Aj4anwSuMJetofwYmeo0QY9YL1CRtcndcth1jWgsMuKG661GntEkO4E/ZRMxyvI9FolNKU7YTbzbf3w5mB1Jtfq1k3tzbbr/dskkW57jBfXkOXgWsMGrZ6gNLJS9sibZvEHt/SsIBmL+bZ3jnzd6pPA06VWlh0dHfkHhHpVr+4zyO9giWhx/e8oMM8qK32ZQ8Eh1i9ikwoMAps5xR5elBHSNhM+qc6IrTkkPOukxq0b7q2ygWRnXJkzFJnotJPK9mVTXgGuVt1HuS70pwFZrLhg3Qu+kvEhxiFY6BD4wR5+y9TQGi8zLKoCnuWhZbanuEIP0sh+KTvUjzGTgmS8Oq/7ruZ/Y63rjFK7fltQVg1Fu+lFnQTdrE6MIoBwr3MfdBQIo4zsKhieOtccubqVijvjRXI/d0I1Iw91211zheAytNbrq2qTDco+9WOLarYb8KyYI2clHuPb/4hjeeAlPp6j/pwHMmnOahAFL7a6p+jvib7OeajXi79+7979r4uX7iotEeVjFD0OaRz5XbQAd46RhgWGBYYFhgWGBYYFhgWGBZoF/FD+OWvgoujhXi7vjlY7/M5v/p3p8vTkE3mh39dqCIJkLDnRx+r0GXk9YCu/4dWXOeG8tmASD+qbD+G0cSQFBrgeNnXywKe/77tdXvil/ao5aKmHVnLkoJx6ykiI49PjUbaucjjZmJwEDE5L3Ejib6EVXPZEwvnlwMmjHZj0834RNAJDOTZ97bXXpuPDIwdqLhQgw3GKU2fnC7tJWGiRQptywVYbNGd+6otTB1yPQ71P0Iisad/UD3zovyr1sMCk3ufBhQ4p8gBT5duU3S6nk9TrSD10sVHwaSfFXpQjLvQJsgQvvMkjL+U+ARsHO3jkHD1+8NLWw0CP9oIp+rE1Qdjf+s7vKui1q8BCYEoC20p8xAwCKKVXods6gMhJwAgFm5Je9eXgBtd12Q1/3Ck4VGKU0CdnvgkmegYHmr1etPPhiDceaJUUgQYFCKJf6cg8quAMsOmrwEbVTUN0+1Vf4RH4zdzXjPixRx/XFnUCSWUnXZfSgbmesQefzc25TinnmkvufsmQsUQmUvj2ZdqS0t/n9MGb1aB85RaarCY7PT0V3+Kt25MT8oKLHFz76AI8+POeVypnpRLw6Oy9CbWaCJzwBm85WOFUQc30l400Po0nAtC3mYdG7m3ceTJH6dtM0YF24Ei0oQt53085NIp13T9oQ5bkJqITK6YIumEL+tiXK3DZOD/6hS647CO2q+BR5HFbx4M6fcTXnKuc+RJY6KUvedrIcwBPSp2c8UUuXgHnIFW97BKZsUcF30r3zJusRKROMk3BMoau+6cJF30Sna2Mr8pszv+No3v3WEHmd37bjPXfbmiNdLctMFaQ3e3xH9oPCwwLDAsMCwwL3GkLLK5cmWGzvhhHD+r4tqxf0MqW//Kv/pXp1371V1/+Z3/5r35Xr7p8T3Cvy/V5Tb9Og3zMnwAAIABJREFUg8Jm/Ty04xPL9WYD43JwrtXvB3D12wng1345K/zOTXv4+4d/EeJZPc6CyKoFh6DhShrgwGMtBf21YkzFOPxup14JWsDj0PTOWPUuq7qkgeHsoDRc8HKwNw9OqTi6l1ULl22FAjAk85KA8GI1GPsXUSZdg9u+PmkeeObymq7syFOuQEIcHnLgeDULuqxyOT4+no6P7k9b9yqQ43brtQR2omPv8tgxVYN1sTStLLmjb3SgmzK0OWxv5CfYofbZjlLLuO2VqNqLRzZq9gEX+NCnHtqhTx8OX3ilPbkR2qle0SqtmF9eKSGZeIWQr8RlVVH2DqpVNsAXLK9gkSyFiuwLBP8trZzxuPJVU8ZIbR4zbKB/CQpEfoUvBC+ejJfxFbxoc0uI5lGyVJl5wCqy2AMAxhYagNPOa3xeeQhPCYhN9hUMfXZSr1jyjU7gEZ4VKC5Tl61tVs1FkgNgLFXSmCxJMDjRDGRwVbzhy46FRqXALWv2BGsRmxDCTpD2JlEg1vW3o0CFx1hVj6OEvFZg6p233/JrcFqgpQ7kaSuGZLcEyLCvtDcHVmwhBbqJgnBauckGbfMxdPGiSHsFXiroUGNasxBae7zmKcEpu4+FPaFpXYqgel240UoyUmAYbxJrYSthc8ndaDjCZpgWfLLgwtfcAAa+PjQHuIfkfkDAA3kurvSVS1Hfm2EreOiVcWLNVw39WqlMbnrwrf8SpwaQlUbwiFyZX+Two4+5TdrWPAAO3vShHfUdrmONjYDVB6DgVPAuVcwLcODdEmXmPTFY6Of6q3l8+5rGhvDjT4VQDG8dRGOWu83hut6Qg3ut+sWPVVICRNDp6rxeKQQvuOghq1mPyEdfn5iCHOw3x6umJL9y2sB2PUfVpmWP4HLfDQ1rLXmYreCUTSN7cQE28CmjM3eQsk3dL2kjQau+Jiu6jE2zBbRJfAWVVzl39/Q3xDExxmLRMWMNvPmAL16sNlOfbhOC1s2N17K11Htfg/fO5dXFV3Vf1JcjoFVwvCtao7pxvVuKcborFqhZd1e0HXoOCwwLDAsMCwwLDAsMC/wIFuDh+xWJp3m9zXilvYWm6bd/6+++/MEH7/3O3v7O7+i5/MSOVf2iTYDMQbI8rJPHGYAusElxAqjDNw/71Be45kh0eAt8AkLLY13welqv4l9tclwa3U2Y4OPaeEWWmCIvRwVfFj0SxBIx6wEMwQ106nWE5iYfYAJXtFVv+uPwhzYrJijjULPh965W8+0f1tfxim4F0iJ3b8+eJ+2pA0tKnXLaevy+PfSDQx1YDuTv6+ABF5rUgevTF+H1MD1+2sGjHfpZRRPewPR8enzKHBmXwl+cWvrSBp1N+UM7dJgbGTecesqhHRmApZwVI9BY6RWxK+0pBn3mGAl8vNR6ja0CF2s5zafasurZifab08W3aqsxI+eNVmGxB5IYiG8CaCLSghyWQfyl9Gwnrhb4QCOpZOVaK9g1q0AlG3SdWhnd/CpXN4x5XWwOBikwZvoKqD947Z7gKygWO8CL/ZSSaI8+3iftc3LVePZw/bhwnXCQQie0Mx4ERvdlP15/Pjo6mA73D6Z7R8fTgV5j3d/f9XWVa7ZsUTzhQ0KftIc29bSlHBmBoZz+4NBGghfXMfJwP+HV6YsLzQnZHZ7gBTY000edOcMBHDr2/Huenl+iFxvlfsKKtRrS5b4LHQJePa3wTk5wq2xS91yCVnmNHb3CG/gkynxYBN4VHFuCOYEJXl8PT/ooB4Yy9lrGtlYEph8alKWOU+yZoFZoJQe24Ou+ndV9fuVWfaTAMPehk7o7derHIH3kZauyGeX+nk7d4yEWlJEnifnBAd2UmcPQpC0JHHA5uIOQgIEuRdtcn8NUTppOzk6/olXIb//xP/Fzx450C0j0MHB3RYM60l20wFhBdhdHfeg8LDAsMCwwLDAsMCzwD7WAnpT1gK0H9vlZ3Q/d8mBZ8rHSghk5yFfTyw/ef+87f+Cnfvrvy8l7rh1+vsYv1FrGcy1nHV/Szj6MeOr2gz9EW5kHeK+8kbPBj+ak2UFQXxwX2hd8HAjRaghyt9LZnu3BU5OciKxwkOsJCf2avrRFLV6zYdUKbgX773gFmlSMmzCvSGtye0NwaeZghHAwB46/QgGiYyejHBfZoV7jwrERjxJBCOIjWtpFZjrDUWzBLwyA7ZAhr5IRcKgkR5L9qPRLP2nNKpLdKzv49187llNfUHWGka1lOeqLoHKmmvxxvmLb5OAiF6lvYzw8TurCfyoJBCvRAAeWYIZXlqmBOmn+Yhx2kB6ybPXZ0EJsuNAOTs/XNJo8KQf2VXC0eVVZw6nZB6aXW1CwHEiiQdO5BTmFp1ko2yI341/OrFepAEozNN1f+kILMmUX9VEFUHC0eXWO9E6irxxXACtAwHistVroyaef+jWxN7/yFQdndrWSg1dv+cADAT9ew9tVEGdbq4J+67ffnU4vtLLtmEUf8HUoTaJUgDgBCgc3cKJZqYbseoXrZq0B83xqDrjaPbaiIQDrg7zMMW84TgQD3LoyULAOtwGp5LLsjjHajcJ7LMnkN3qtUgAlm2i8rleCdzR/+KqqrwsmEJgKtgtbjjyR9yab6kwozxuWJLVkG6fcrgVgvJrxGnriKBroRbvrkpFyVmvBi+txX3b1GKsOXVYIETjIWF3pVWnzk1517XCR1VgzFTK/IxN0ObATbbWisco0kyKT5WONE/cRgiySb3eLVy13FBi70OuR55KFAB5vwilQqgsc3JmX6F+yV5oCJ04Wq3Rm2pkPcqhTWZOnZOfLiMx3VvJCLzItc5k5DC3Bi6f3JIOJxqHmttbOmbb6Je/aNzZwKtglJNOlueRFCs113yexB2OtlWxq9fzT+ADH8EE/iXs2/dBxO3BlYfHnNVOtVpNMvCpfgSPBM3clEzrlww112TLSIqRVzNAKX8rw5hpjnpu9BLHc0p+cj8rQLpIlj/7ugWceLVAlTYVftNHAdJWbzmaOAdA3c112EefC96rl4s/lTStpj73HVCFQx8HqZlbo2j6iBZ8Ehguj7FAyIVvNCcEpceHAY2v77Xe++sav/er/du8v/id/cfqP/8J/2KyLmYUDw1zTwreGzV4mOE5fagtwfY40LDAsMCwwLDAsMCwwLDAs8I+2gJ+25TRpr7ELeWer9U/99E+8qxUZvyu34UMcgzhUPInrWAJAok2dlLwv05b23mkzQsOhH6fg1XgV8Eh/nAdg5fba2Qh9E9AJeQ3fXqcpx2GRMTTAA5aU8i1acrhZGaEf6EWv8IHHsY0Ta9s0GugXJzF0I3fgoF/8m4yNN44Qr2Hla2XQIgjWy4qc0LklY8PfbOth+z7KHJEPuAQQsCcpMlMOXHBehf9FcJuy9jTACS3ynoYr7QSNHGkPXurkacNuBDZfpUN0CR44pi32mzKEHkEDBw6Upy3y9Dl92PH8/HT64Yc/mH7w3rvT97/7D6YP3n93evbkyXR2fuKgMc6pAzGZM4rPfPDx42kLZ55gTpMFerxGNSemacMhcKZRqrrgnFpGaI0E/pK6a4t2DuYzuWQ23Wbn2M22Ciz0CGqovq25X4E77LGeDo/0CU7RIpBKCj4BPOATQOZ6Mc0OJvCGE2xwae/bKJN4HS02r2tQq8a01xdlAmN7LeDEq2q8UMZKPfgCU8GW22XmiunZFMv4hl9kMHOdgO37+nrkCg63M/ShDp/sS0adPcnYm4z5QqI/R+4rwPU06Q9tcpL5E3HRfY7N3ZNo534FGLCxK2UCmfAlWE89PIwrHLU6sEMfi47Ik8zP7WUr6EDb9FSmn9TnoZ+29HMNQDuy0Z/6+fmlV9phC/ROIJEycOQzHRWpZ3yTZ34YUCfaGQNWaYEe2vSHbtEuuYKXvtSTR1bkz+EvUzadsF107G1IQG9H+6k5ONbkQBZ4xwbkJPDSFr7Jw7/BqepEjE2v818/0AdmX/+lX/olddtm3ADmgQx9cL+IPn0jffks0P1F+fIpNzQaFhgWGBYYFhgWGBYYFvj9WAC/uB6Q87xczrNpqUO/1Gv7lsvV++9+b/rJP/hPfXB6fv6u+p7r8fvBzfpGW9jIw1Dii4Zq81P3jhxXvtYFXQ7a+UHceer+dVuItOsfzgMJpyJOSOBxOFhJQIIZdZwar8zA8TBNdxug6vCFdu/4qRsfVLSAYZMW76JsqZuzpbL5t8BCo+rgG44fMpHA52AFxq70TYoThCDABp4VbLtyfOQ+ocDsRNEPXSc5tnopxzg4pgQaBKpjpdfF9tReNgS2dCyHqezjYbCciF5S3obr8SIXZkh70Skc5C8e2L6AGAECNtSliuTRODCO/ENx+DKhlJA1eNDF6YNn2sLfwDrVmNbqFOxPKpiiR/0WrmSg7jWB4ssIFP3GP2PMyhNPFvULOisFw584ArxrvywR8ZIO9NUIKKMEbNHWeDe+anZCBvrQDzpwT/CIa+Dli2fTkyefTVerS68GefzoEwdDvvGNbxr/ePe+bNrGEYZS/emz5+LNq2y1WojN+tftS4YWCKGscdlJApgWGno1GfSkc8ktO+kfY+RE5ErqOjFWM65ouV3QtLMassnFVyJvuMxFE0qkG5YCMT9Fj69lXq+upn3B8Poi16XtAd5MX0is0lGdDdZRlHHGZr6ukNCwJRzjhG2BpJ0hqglWgRf2aSIxtPDiYGxq7iCjjTTrYGApCH/oAu8kwqzWuWkRPXWVHJCAr7JaJdbkUt3zxcjpq3sGTdDuDxRALX9pE+KJHLICSjbeU1sFlG40Ly6mo3sV5FNIy3y3r+vVVGxwy5bYVrIz4/o+r6FCBvGBr293qteefWUT5JNERb/ZqdqQVTZkHso8aUNfRp4EvypULi51/9J1A3zJQpy17Mw3j0ms4yMhEySYYrUardmQ1WyMg3jPK2uhJ868asr902OsASfYKdN57MXV9PJ6ZPtzJBj6Mx/gK0rQYO6xuMr8BSMeyI3dVBOcLIat9U/NnBHbcC5YAaO36x34ulbA9xeJZS/4lT10h0IWI4u1/vnvi9pSxrbVVvPI96TG2aKaJ+O5HPPfQ9FhtWBeYebaE62tWmnGHNLf5a2Do7OLyzcfffbpscQ4Vb8W+hUtrgfoknxuZTeM05feAiNA9qUf4qHgsMCwwLDAsMCwwLDA78cCeUDexK12vVyzsz/977/2v07/3D//c08uL1ffPzi8/4FcnsOrm9U+DhgOlB72eb6WX17OQh7mqb8qhSdOAinOWJ7P0x9nNM4X7la9CtUe8OX09AnnqmgV3fRZRnk8/GJPok7ApLkFxgEvfHg9y7LJyVpkKcePOnoBS3AMx40VCqTAhg51Dl4Tgmcck8CJkmiBW1+hw1kGd34lU54k9Pla3c5OOaPgQif8zEu0SZRJwEQGcnhvjkX1Fx52qLEr+zXyMy0XdApNFaos+cyr2Yl+Ujm/oq1qcGadO+JpC0yfQ2dTZtr6RLzBr6/N86h6Q7fmSrWVE7xgF0yTX83hDQQBP2Z05g19bu9kd0M7xb7MP9uxzQ/2Trp//77nHa/Sffr4sb/2yHyJjATwWGEFHvvHP3ry1K9bXhPEkX3X19ofjDmyyVt10xCcA2IRiPY2Hwjx0GfdrIDGBDoc6ESf2hPYxEuuzf0lD/pr3hoOXMaYunBtD+E7GIhTrjJz14EKB2dKNnTyvC/3u/CgpYTsHL3dq6fOZfPq51qMvaBJHznBNsqsGKskoQWbwALBCY/NBh+0vhE+CXwH6V4hT3gasJ2Aj+w2ntpTT+At8wYZnTCyErjuU7tto/EhXa9uvFr04up8Ojw89H5pvD7oOStlmC/gwYecjyTw2uG2ymkH1iuVCDQx/sxh8SNFD+q35Fdf1QXDPUB15mC92ss8avcF5Yw/CVqULIuC5OYrPbAhYMXDoJ/jhc4lS9EqqDrTrv9z4lVirHOhFWTYlaCfVwOqTL3oMIVlS+GlDgHKyMFEsDwKYjkXYIKvxagCsQlyeZ5VxzxOptPRtJytLu7mRUCQD2AkgGgYyXDNTaTZhDZkDT1yz0PLWvJm4V9gmijmEZq0UQYGm3seabyp+/Vz9WsFob9UyRvUWol8vLtz7+vf/OaPf12RxXf1cZCVYD0AouOhDJ+R3y0LjADZ3Rrvoe2wwLDAsMCwwLDAsMArLZCAUjlmrwRZGnnqV1pPf+1//B+mjx8/OfuP/tO/9AM5Z+/rafzHri5X+zhnSorX+IFdP0jXazZ24uTEVNxMD/R4qnKl8tUz+nlGz6uK2evLT+uiRapn+HJA+GFfT/12AOCYr7PBl2QHSQ4cbMpJqEAFX5T0SjPBkOMWuF9+Ae6J3QP1OXff4sTY8ZB3gxNSm1yLszxAggCsXKIfx5XNt5HDsrRAEb5kbLC1pVVhtIuP5QO/wYMDHIcDIcCo7FU7CkYQKKPOq3orrUJCFmlrfBVk3hpHbNV8HsM39wcIwNwXW72qHvnBg18CXEUHjkXDWjQ7mZ867FRaDHiV42Y8j03JBX3gIwM59utT+pPTH4cPUgVfdo683shafdkrCnqmjcS0WyThqD10yUnk1xqQBM4smxxqw97ggAtIE4t2zyFk1mbz7leX4SGkhGzYTQPX2mvVXPHamg7v3Zve+epX9TrdmZ175kwSMLvbet1LqwRZmPVcMOxN5kuGQC2CKGoBX58igPDM14KKt+o4/9Zfc6yGpHR15IK5c9vkxqlgiuDoR1euW83z0kfMRNcJ/Uipuyx4YPX67x54LaFTbx+DNjzavVJHjdi1lCp4Ah81/4pnrk/NBI+xNpgyB5lFdtTIye41L9ysEFEpqN0TbSpowY/5zLXDdbgtec2Xec6Fqn6FXMwXLPPXrCj5wQekyUOlS4uO3GeWjuiffoI7JHEWT8ncgOtDC9iDr6nCh1cuz6eXL0+lF/tS7TtnBZiDQg7w1JwFljYAoElyyCVlVqnJvpEhlq693LBB8QMPuyhUNAd4at4CIzsgu+zJ7wltBnhOco/SJpTCbsEZ4aNhjV/RhirXcO7vBIwI7mcFFLO05OBaLz7cs8Pn0h8yUBBIH1fgXssPF4w3cvXjjg7U5/sFlkb2ZiOmGXx49ZQ2/n6kH1xJVWcDqq6AZRJzwv+RuzVmXtWKsdK17Fz38uDmQxqQ9d8sCiLG9W547E5UjH6VS0aNpeYoiesEuPAre0v3dp2r4L9d0qbBG08VWRx9oXG9dXRyfv7tg+PXvqUb2Cei/QLKAlA3vFFsmScmNE53wgIjQHYnhnkoOSwwLDAsMCwwLDAs8I/RAuWn6PmZd1b+1m/8TT1nn37ntf2j7+zvH/2Mftl/oPdf1Ffv0cgB1ZtP9Yv87HwIdS43wXgeB87BnvIDDEN3vQIX96g5Tf3DP0/8PP6LBkc5RRBpDgJ9qsVhUBFXgLPhqZPsPSjPii7oWHbBUcYhIQeOvZ+utYqHNhJ8kR34BMdCjz7g2KuMhD4Ew+BzLX8EhxWHK/BsRF1Bxfoqn3EVFIsDDRy8ONiPrGRoRmuyzLRw+PGKzJfgD8592Zp2yulLmRw9sV/aqANaeXN+O9om0k7Bif3T57FVBRliR2ADH3mKx2IP8MGJHtTBwZcr3MhbY0hbTwMH2XUHQcoW0Kh5RV60w7/6ylbhCf4175KC53PNIRxYt2HjTpe0gc+cIOULhAQ4X7x4MT18+HB6rNVj33//venb3/y2YQge1Dxic/ay96WmzaMnzxQH0ooo5o7wt7R6jPkjw+gQb/jrsA7IpPbYaNN2DuzhbDeH2zTMXSQYZ9F3grb1qqptjQloc0Zgp16lpE4XNoiB2M9pxYcFRJPDARWBeEP+Nt9rPiJ3jXfJXPQhlDHx+Ik0+VrXhxOsJAtt2Dib8VOnneRccKELPw5FnrU+s1Zmsom84z3CKbwFF7o37RVvr5QTTeibhjkUD+gvPMTQKfK36wXbKAFXaZnjkbd1WA7sF3kJBJGoE0+BxCUfE9C9NnzpN+1uTpZt2FeLe3BdF3yUAH6bPBP0IRRFcAwm4jDbJvQdSGy8/NqmaFkGhNJ91VkL0oODDPRbNtUrGLbYmOvTslgvnaoL1AqK8boibXSJF9cHdthTYLr0y+u03LMWGAiZrxCLd+mf6xHcwFcROO7nS7sBJHuNQ+GblmSxvQQQvYA1nO4T9FEm0Z/7hBvaKWOQQH5PhzJBsgqQNfnVBg5y9/fS4BHkdPLQlR3pA0c5FlRcvWyie9G91frgJx4+eOMnD4/v//b582cKkKnveoXyZW7hjnT3LDACZHdvzIfGwwLDAsMCwwLDAsMCcUDm59/2YP1FlrkNj2uAByAvVAGik+cv/5/f+D9/5xf/5V/6TTkE/6IcuW/qlUtA5PXsaOGJHrrlbN141dbiCDm4Ue6PHYg4PuSRhgUKJPY04uEdx1Dddg7sJKiVX+BxAjiWFQAViLqGFq9/ib+dBOEKElJOrI7g13LokggO4Hg4kAYjtdsplg7gZ6UB4MAR6PAqOPtTBEIIBJQDY36SCTj8jMgoKa1D+SvVDqsEK4CjzAoeHCwCZdCgvOJrlugpwVbtS3sEyOjntTI7tuqP/YC1PeXglzylA7pCjzZSZC3Yao+8BmgnRLN8GIYkfL6+yUbnhmfxgbpmug0MUOMRTBE8NqLe800d2D5FTmB7+PAAdpZLMEVH+kk1po35NoIVhEHEpvdsqYIDNvDwLdrIWeNN3TJcK+DVgmqAOf6FEErgl45lk5J5sffZyel0+uLl9MP335+u9KrlY23ODzyvXFbQlTEvWuDu7u9NHz2Zps9enMtrPfQLwATJSn/BIRxGx6XVf89vBGE5FTPFwTO1YnPalZhb7Nfl+Bgnk6jrJ69Pugna0Ut7pxWgSfjESpg1X6wEDkPI4FyX0PD81S3gcPfA1wlzFJkJTnDdXGr/NOoEDa9UZp7zSiSb5aM/feTQy4oZtIMOejnpwoUegTHuGuyTxZhzIL8QOU2XksMBIvRWGytU+w3oPWbiB0/zExzlrPDSGiWPkbdYUx/7/0U+y+HTIjPc6ScvXRClZId+jpVWJPn+5YEgIIIphYcCJN0zGaeyQbVZ39JO7YcVySjoxrN4wY+U6yfzGds/P3/pvnzgQZel7QNtDr7eyOSAL/L4SjC5Zhf1zUEtL2kUOfUvX6ss3gSgwefLrLYDK5NEmplYdsFG4NZ4ykLu12iZnvnL3sByv4QWlK/bXNrbg94iJ3Dc01lJZdistBJ/6y/d2M9ySwOJnosMaFj0kZn5RhJrJ+CS1oyZ2Ca5R/cCr+KyXdBJ8rKSjrqsx+pLYuvZ860fT9tXcF64lfsiOLqXViBScgkXqg5eSxauAWyVHwi2mv0kscdMZ4snyxmx7MGbt/o5RmPqr02vpqPV5dW3ju4dfuv87PQQBhUU1SzURqLCLCNE0ZHfGQuMANmdGeqh6LDAsMCwwLDAsMCwwD8mC+jZmSQvQ9uWTDv7V7/y1//ax3/qT/1rv3t9s/7h/t7uHznDYZWjoadzPXbLwZJTgpPBY7tzPaSTescj5YIrx1JfoxeUvBQ5Yd5oWTTi6OFYJAUHh8COhINm5YDjELi9wQPLv3KgmiqtD8eLlD47aOoLL+dyYoCLvMgDfeqU2SsoDhCOjJ0ZsYncfKwg9CwL8qgfnKTqL+8sePSFx0qbn6fOflbesFqBiMiUPm9Eb8g6QbeHSRdt9MGr5Ei92afph0MGTDOXcT5Ps/SBNnA9P3BTD0/4Rce0BQYa9GNDHNrivchZdro9pyyPTEmAZlcb2RPMgAY0E0wFJgc8wq+nZzoem5pTwCVZTs1mzXfTQS54hGZkDXxy+gmEvfPOO+J57WDQV77ythzovemtt96yHGysXXbT64maK2yj9fH7L6aLS7nEqnMV3eirEqzC4pVLfHmujXnuNl1FDOMVawiaqKqMNXNYwVZvxu0rRu30O9McaeNEcOaGV4E1FeOMG6idoCEDm6ab4ClZFH5wkIw2AuTeTF18cMwZS4IUBHZPTs68kk6OuoMOseGDBw+me3r9lFVTGTtsBy4JtWgnYE2OEVwXD+BIm2PqOeagBfcT2UCiMrsD1+eoAZ20qeY6bT6azcKr5i+2hmjLEUKpYOCUcvGEdvDd2U6e4y0AQ7/rrY96ZCJ3sEdtSekP3Z5H+oDlHnWlZYmReyW7EHDfcdB3pYWKNZf5imJWnYFvGoJJ/A5821804YXdKv+8bpapzBBxb+lCo19thZYDRqU77fwdQEvQ4cn9jlfauc44/MOIIAhAkbjmScgCvPbXck59mSfIXoZOu0Ctb2+r6EOg2eR1SnDQ9FFaib8CBKrgRzvJNtO1QI1ybJU+cv52JGV+AwsdLorCuz2nS6ayCP2Nncm4TyXaSTMtlekTD7S8WW9v7V9cXH3jtXtHP/aL/8q/ev9v/PX/GWGMAqhL43QnLdDFf++k/kPpYYFhgWGBYYFhgWGBYYHfgwV4bp6fnfUcJZdma2v9g3ffm77//Xfv/+t/+s/8oYur9U+srlZHehbXns43/LbOr9YgycNo2HR2D/CU+7p/dRdCbYrfHvL1XM8rhsA5IIXUzTPgF3KTd2CsPeVTFkOOmbGkwH3HUcFZUMl4ODzUa/WAHB03C1KvUeJEEYggCMEv+KTV1fV0oSCV2cvTlj9n5/1w/3A62FegSv+8SkaOP04PtEm8MrWr1+QINlxq5c3Tp8+mc+0thGN33wEBOVNyjHBY2YD/Sq+n4biy2sUOk+RdKxhwdXUpnoITfcp/8Kd/ajo+1moSOYJ2/hUAQUdgOLyfjSWoU+RJEzYt/eNUYdqS+da4YD/BJgXGkF27hJWdGQd6ytkzHo6vWuIUgp9j03kEHp3J6QvfKkeOcg61UFF0Ga/SgxVtfh3VclgE4YuXRAIfv5g55nmmIc3ePTjb0UlYc9mmYIUWB5xmXauNLw+q0fKavniEVuknnZkk4shG6sfH96c333hjevMgEv/AAAAgAElEQVTNt/ya5cPX3/DcYD5CGvq8Bnd4Txuzv3E8/Y1f/3+n/+PvfGda7x9Nq462Li+RxNaRVfgoR/RHibJX6ymwJmVg3xIY6vd5bnS/9S+CqnceMzt7M79IzQ6amCqDr3aNAcJ7M39TVpvm/v7N+fRv/Mmfnd44VtBMATVWl/mQPS41f19/8HD69re+Ob3z9lemr7z1pq6D4+nk5Yvp9ORkOjzY19xV4EPy11wgYKA3TaWXN+K3Qtq7SdcT4+3Nz5n7TTMUcjADmcUvY6tSUx7ZOWpMsbvHFj1sLyjVNb+MOXEL5glEuY+QC14BFFvLZmj4TT6v3qOdgKZygjvQzxxxkEfj6kW3yOBxFaBgdHaCPziWUTrSkbpfCQeqhGlca67TLAv6TDf6QNWv58LLU7f05ou6To0/8A7C/X/svXmwfdl133XfPPx+v56kbk22JFd5oIAMEHBRUBgSEhIClfxD8Q+Dq+xUKlAEqpICDDgxJnaFOGRQhbhwjAHjYIeYpLBNpLItyciSLUuWbcmWLTmybKu7ZbXUre7+zW9+fD7ftde9573+SY6RWsDrs987d09rr2nvc+5Z666zD7y5piIqY/OYnjj489okjEvBJW6bk5THBuWRP5dNn2Pyz6jgE5pq1mjWLA6mdsRO9S1ezyvTGevw5s2b+W7Q0Rfd6SSzH8Ael/UiPGsw5x44lEd+yHLkRxcY8Po4VJfx8uDRyb0mdcqJU2ebqXFknVBXr8vvJXDaL466Hkij8IU/ytUvJvnCcSUDLiCnlrI8KZvwsuLaaAe/oPWCF2Sh3OvAPd2cW8d0WwiA02Y6nBf3PODXLeLaNtZ3+bHl6T/+x/7Y+5999tmnP/yhDzoNBBCJldPJcXN6xWlgtfJfcaLPAs8amDUwa2DWwKyBWQOzBr5gDWB/cuOOwfOB97/31t3bN5/e3d76JJEfh9yke5/lAQhmE4c37R6mzlMZ9e4f9v0wSGqccI2jx8TYeEl73d4V/mZBY6Xu9s0bjzApY4z40IopcBpqGJVtoGjk2O6h46sfGRK+cZUhVNFOwrRjrGkErwM0o6Brv2N9Qkk6JnHEyBk6qr3I4FHHArDiNReXOIS3bhSZ9X5USVzW03apbF/LYvlzpeZ3iqNhp+Mv91uvR4MK2seVGtc0v1xuPI6y7KF8XVfOLjt2Cm+7bR7RIQZ+cDjlOhNieQq1wm1Z2Oajxq3WQONvWg13GYdwzqXHlN/peMdMk5FR27v7iSDb4BHK5sP29OFIdU0YfYXPdfHMp59dHCsTq1JYo8colp8K+TSeTeW4QQY9ChMdxT2N/jTS1QaLJoc8Klcfnsvpsx36zMI4KxgDXA76lrm4TGOeSv4xN8NZIQ0f2cs5LV8kI5N2doiae/SxxUMPXwcd9FgnOoqv8VbPR3Ee6vxwzsXZ0UI6xXQy+yZH8aoj+4uubEW6mntlmMqGjsTXh3z0HFnuZJsw3dd54za3v1Pwlc+EprreXB7T9R5jfYqn6dnesJ33GPOWs9usT+HE2fXm13of+QGAy7JrdQrb8qzGej2qc89rij6hErnoxX824dXHC7MxPaul9hcrDpsH86mM9jbNhmnZ5KF5W/G9kquvm54nwvW1U5xLfbjYOKTh4ZiWbZwqtHHe8rik7dN+8ZiaH+UuPPUjSPNk3jKoqy5P+y/LJs5uKyq1BnWONQ/iaThxNXzLZn/D2m9qmt1+mZeGCTDg9KMGZUem88VjW7u7j/zhf+2P0uP5o/JW190xZs5eQRoYZ/4rSOJZ1FkDswZmDcwamDUwa2DWwBdHA8Oaxgjh7/bN5w5uPf/ck3u7208S+XEfW6CNDLZjGfEz3IBXlFbd2HtD3zf85t7om3vznht4DWfwWEt0iMYdRnbDmWtAXBgbPN7oM1CDnEOjraIsHG8TfCSqYji+gMEdAd6ydMUZw4R8HWO8jJSLxmhUaD9Guv0xYOD3hMd7lNb9wuTLZBSP0XBtzIV/DRTat3lz4RoRMmsY/0JHfsYZlRG+Bw73tGEDZSJ0Cmd4xI51w3KjG8SZpDMCfpo2SPJIFBSqn09h25i6ADsgClWMJVpW40AL7hovaHigoeGX84HuT9Fx7RskZXQH281j6A9Lteeu8U1z4Rqn7Z1qNYm/IlA06Rp3w9QjvlWrNVd6cZ5M8m7KOOispKy2NlLlT9jGb750BiBT60BcLcsU3nZ6WAOF1/EegTHyMVEzUGfe8GBR1TFFomuwurjjixh4wx2LkT4RubbluMYHkLGeMyZxQyTl1YdrQsfIpEW9ua40lzMfjrGxeMRLRh2eHMMR3YEATDSUXigUo7aDY8PJ8BE3cBi94yOlOubO2cPMcZs4/YQxCoxgFrGn7rmhcziRNKDc2WU/MpwgmQc8fIiXw/3GjBjbxsmWlRV2y5na9ZJxyAAuHX8Rm3NB9mp+lME1AQdDXnPTNI8uacv5RDxsv2hAmDiDkM2IKGNl8/bY6HilZMfLl2/1dIz1xtl0mmavzbpW2Xox9fiX9Ms3h+d045bfunSgOFL4NXIrc7e+OMYzcs78ep5mjsmjJdcfTR7WG584inevk8juOmG811LdrjlQbkf5Ci9cjuCqsnz1tUc5Eh078qblmJThRR5KFnTPuvea4ptdjcR0Dzx57+8Uf7g44RqOaKw9eIRW82Bf14+4Nvu474nXaeGUxfNvJGk7Tv3Ja/0w4Y8eykAfayZ8wZu08p1E2VPIo/UoOnEJk+0CVCqHy8j98qJk8dkfPPUDSK79EEd8pQchdDlPp7oLf/DdvHtNKp6BH6nltd21Zd3D01GQ0X4D+V51cnKGKz78wj7B3wBdTj0/l9vn+tXSwEtn/mrJN0sza2DWwKyBWQOzBmYNzBp4uTTgTbaxBdxpk52f3X72M8/88vbm+oeJfOGVe/TUXjCn3JxzL14GUhsfOnWmqW++k2s8kLyZT57PqjcemywL0zitT8uXYXuMuQaFxjjmQvAIa3K8hwa7EVxdN5dWOX4KtvELa2SLyTaNKpPwLUPjrHaNLfZdwgiJETScG8JkvFYWqXGZN32deOJv3BpvrcuOgrOvjW3HejS+zu0X5zQ1bNPqfvPuuwyvCdep4cybvn1THWQjaNqafuc9dorLtgcl2/uwfypfxsTorLmNH2kgEa55selBOLq98+bPeutgJdtqnqY8NI3wwrim4zrxmOKyHCOXdci0hT9xSWNjCycAy+rXn3wqBnztyXdp3sbcQiSYltF7tg95z9xIfyR5Kx2NdeFaG7DBIZ6hd6N06MRJDU341oE1TZGLvjBOh7jDu2sCvPgRFnv7O4sb+/s4t3QU6RgoukaBOb74SU/WtWv5+OSQN2mWs8fHZU09D63LzjvqTphus2zqObHcfeblDKz+nquG9xwSptMURxyTOidJU3w9p90eAD56rHnDT2GmdGxveMvTZPv0sK9xWm7cOh1bnimuLgtn2VVruedLHCbr3SZcwY5znxPJiKtce4Zjxv7MC9evPidqnlyjKz01rqYvLcuXU+h5EpB6TMP4CCtOnDirEkXIeuw1IcwUnzI4j7412MO3fU5lq3JdCyRnhFxfs8XVtIU7XkYDF7/No30NO83lo/my3Hx1nkF8NB4dd9Jumg2Xx3Gdqwmd4rvgu9zjxNt0Ldve9C1Lo/sZu+Z4dYTs19c3tt7wZV/+xtevbW5vAOvFghCzyHdhksQzp6uvgTpzr76cs4SzBmYNzBqYNTBrYNbArIEvtga8g/aOWeuW0Jbze7/56x//pRvX9z6Ew+y5bR6h8iYchw6W1um5kSPesHujnl/zufX2Bj2GDEbCMXfq2F/Lxxe12/sXdn9xP3cPJFJu+nEm2KdjwaNv3LseQD70s5WvTYOtIh+ah/AmDxDSieIhHts9TBt4JzTrY5yx79gRPPjGPbsxDYl84TGfYTDrqNJ+SPQYMrbRA+UYJhry4pd+ElEBiYQhGmKbY9M3Ak7GabRJR150Gpi388OyDjYjdDSKD+7dL5x86vRLgJEISBpFOqXUM7UczcM0l7fmz/bLfeJZJY1ma2U8N2zjkL+UnW8BmXu0Fh5sz0gyyyVX4bG9+23v+ey2KV8Na5+P5jV31l0VJtuIhUj0hVEYLcOUX+kkxI4oJVdU3og45G+6q3UUtHnkVXzlZMX4Zh5USFQ+1kP4B7e0jDoJN8xDy5D2EYlSnDJ3yszhOrBta2tncecub7B8/vkl75FPFRo9U6EoNVfKEVql33AKT8vcKBTr6qfbkTfRi0iuPMs04ORlnXXrOdB8C+N4I7GiO+rqtfZYqllI+1gvj7/q1bydkvE4KVr/rsW7d+7nXDq8f39x7969bNp/QH7k48I4x3Q65dFLHGmeO3Euwkn2GwO3uBpfR7/JdkUXqorSdcsqT5aLZ9+s6CqpSEcvLR5xfrte+gDGMUscWVmrczhn8qTfKKS63hR9ddU6smxqHhpv47ZPfMFphTTtU9aWySit7LnmnE+S50vWFUwkgtI55bBdvnp8YIZ+uiwmnaDmnrMeRlkdsxaNuBJHRVJRMop1rCfXanQL/rwV0/XPoQ6XOXqWn9ZFZAS/F12vn32ov3IM1TmTaD/AgmfoWRw6yEofdsIPPxoEt9GQTGTz1N8vnn9hmfPtGL67/5i3LVuuPdQY53cBVylTYKCpio0cc19II8X4X86LUWoq1u8uxTVN5xUXL9jsKOd3nGHqETpdlk54WDrilMm5GusMnfRLB/wekBd5SiQbRPM9Acud99pVZ563tve5MvS/Bg7faFnfa+fne/cPT994597BG9k/cN91QpJ4Lp+pjQ/Xypyuvgb8WWROswZmDcwamDUwa2DWwKyBWQP/zzXgjfT6+tbWyTvf/uP3/8Af+iO/tljb+q2tjY3ft82jgxhXBJ7UnbXGw7hJj7HWxsSKtOaZxlHBaRg3/BTWsih9dNGkgZEoDtoydvT3DX3DWxdfjcU4ZpxljQJhtGWMcJkao+KPMUF7PWJDrnFBPUePHXBt8NgXQ3YY8tLxsD9RMhg7miC7W9vYMsW3Y7RLNEQbT/Gi862iJ+RFWd3gvJwIGGjgcqzGoill6vbnETp5pF2Ds2jQQGpdyNc0tbzTNstFw1I5/YQzrdqHUZfWaXsZaTovom946zHK9yA+Agceczenbp6a18JT/VVezVvj7nbZmZa7v9vNbXO+ki7pCW5DvzdXb/i1fvcE4wrnWBNDL9J0Hi+npm9/4zI6R124tlwXrDCcU9uL+4eLxc1bdxaLa9dDQ14AZNGX7ns8AiIE65m+4PfccNKF8/lEkvhNLpWC0WlMQ6x+8iG+MKael3ZABZ904DHjKCrDGevVlLI5DtFzXmIhvUceeWixg4MMTwvGus6AcmAc4zC7f+te9s+7c/fW4j6OMh0fHl43Xv3E49mjTZzikd9+nNm21qF9Pjrayb5Ozb/14JBvutXxg5I6d7SPRDp2SXepN3ulXfSaB/MpT90+xSE9dRZ5xnq2zeQayfWLcuQBUByNV5iuT9umNIUxpa2KGZO2cZ2Un9TRkXDLtXIJXj0ErjKuT7xUBGcS0wpOHC+s+00cl61f4T0VfGRyqrPmmZ5BoeTwpRb2qUv56NTwXgOnskmneB/rgB8FpGPizKw8zi1qoKuXQMAVNDJu0Cgc6rhoSkMnl7i8tq/7mKyPnbKeqGWsTjNPSGY9cNHbwFcylM4LV3235BHY6KLWacMVHa/ltV5aLseazHSM9VoQLnLSccr5YrKtx6dhfIij2zt3XYWvybwDLjHeA1Dzh6j7oPwK6m/e2N79yOnh7dt5wYIKUL2TJN45XX0NzA6yqz/Hs4SzBmYNzBqYNTBrYNbAl0ID3Gm/510/sfiT3/gNL3z3937fr2F4PLW3s/v6xfnh1in2hU4c3gjpBsHYZe2cqqiuYevkBl9WvREXpm/0NYLyFskYp3WTnpt1rKHAYDD56752TwwFch0J7vtjXVwaI3kbpVaISXjGCZkmjSP+Ntk0XQqaSBoK/tLfRrW0xOOjPpaDFzj/NKo0tjrKwr7Qxth3U3IjvYzI0FbRGNMQ28IB0saxBqb2RxtN5qbIB4Nt7LQsRhednBwttojUg3rxkxGM0eHBmMJRxl11Nc7iTWPM1DQK5kH10iuf4RGIgbtg86ZEmae/YIqO5cxH+qgteaqydJPQc0rUAz+maLBHX7ULmzGYbsZ6CNtJvdjXONPHnMRJqaNQWvZnAOPG2IY3N6JInnU0Oa4fKdQ4Lb0PI1UPlpBa4wMu9Bwqnswv48f6S6RXMNc4x9bcuOJWc9tzDJY4inRCvPjscZyh69eRj3FxeoZXKuRZ9DrGdDqcDocXfCxTCVxV+JG/liu6dp1FF+iYYtbOcKjZHJhMBJyiY1pwfh2MMcIzD1lvOG6JhDSY9JQ3qxp5ts7TWq95nDd0cpopW2hDX5zb20SF3dhfbG6xn9jedukXR5t9knHvsh325zNFnDCTKnhqfQlbzjF4UhfO4FgHGTfmyVkvucWlwxXHexwqzKcyMu/212yo/eLR8z7yD56dAedNyAyEXtEJh8uyy0J88uL4TjreGBzaPU44Ha9ej1x+xccYwdjUL+eApp15yjpa0nB+SGPdyYc8qHuT06hMkOR6VLx5XV6l4tW3KJo6Gg8qcU7qeKIVKfyxoOZJOK8wyQfO6RxUua6XwpQ+S29efuNs1OmGDIkkE0gHKzzIRXEinG3144BrPVPrtZk/HVJi9A2/rseMpc3rrNwNf1hoqC/cawDnCpK2E5zTvgDilHc7iq8fVc1cg0daOul9E6eStl4ohpb7sCWFKdq47ijP6nx2jBFodc2q8fBHZF6lavf88vx2nvqtl8UD3zl+vyir13qEjR4ZrKytb3Phu166BpkyjDUCPMWkzCTfV7tbx2tveOzhR74MZ+AuFxLA4R+RGVkTNbics1eGBmYH2StjnmcpZw3MGpg1MGtg1sCsgZdPA95EY6dqFKwvPv6xj978hx/5lZ/76n/8d38Fj3hcP9o4efQIRw635Nx/50adfU7KIJAl2rkhX92He8OfTb3JTdaBilEZp8W42W8joPobD+bN6HesBq8pRoZF+mI00p5xgQ1I+NiIw6xwyZdGiemUPZzaKabRUw6uNaLjyrgUV2ggRvNjLo8eGj32mxo28MB0tED64XEZDZZoBiSIftRt4StHQ4TRGQc6No0pxwKQQGnERuySke3fQlc8yl/40nThQ76myXrBXsyFuQhb8zMdG1owoUw6Amtbm4Kwb6qLtMKa7ZEKusEov6TmIZVJ/UI7sPLUayK4HD9kUmfLPubDVNgLf+qBT1ccQZGR8SVD4ffxpdANh+JoLKWT1kvTEpttRtw4bpqEcUmI383Gm0dhGtTl+Ozzn42Vuomj1RUkvuhP2RqQvGiXzJ6HF2ezKOdRUIvqgPGRBxmicfEpjzhTpohnYUmLXmksHYfARU74j4wMCyxjbD9lTW4h9/Vr+3EMiNP+4KB/Z3sbx9h1ucnjfNGPCkm6aOTbFBrgM9fp0W0pjI/LOu6+GlM1y6II7FDStF+orju/ljvPWORUuU0rbeHJcYMGAOpAJ8wS13KOVk7O7oseM7jkE7d9wTH4aXrp4zoan8yA0fFSOOALHmRDXetISj7wBQf8GwnmI5TdV1xP5Ka/eWu6wnpd9s2qlj1qk/ziWfrhDbyOnZbhRilod+nV2ux+aVuuenHi+CV93Fk8AJv+qTPPfq/lJh1OcR6pF+o9XpymxmUufVxM5f1RR6HNDyxxpumAU76KyFXHXp/VVeNkwBJn8byS1brncf/wgGSjPs5PHIHS7u+75kvdOLZ1OL6G0iaMOOuHl5LF83uahJnyYrmT87TJOmj+oeH+YzxNu8Hl4BRM67uHh4evu/7wQ6/7d/69r9//29/z3fABj8CAY4WoEc75ldfAxdV15cWdBZw1MGtg1sCsgVkDswZmDXzRNaCZjyeJ90yes0fK4d0X3vXOd7yPx6Tej2PgBQ0MIwy4aceO466bm/c2DFY38t6SeRPv/Xg5DmrPmpWxow/Nm33HnvELt4eG4epXeYydUIKaeITHWvLIW8aoZ+zAIYiGSre5Z0vTrmgFHl08Yv+dQzfBx0BhD7JjIseOLPPL/zFOs0SMpQ9ejCoDtxKIU7n7MIShjdWlAww4HydTB8YG+JZOI5WMiMljkUY4DF613Ty6jo3XCWPnfHHnzh3xQN6oCAAndo3GlUme+ExZmsKaeg7M++j2GhOwMb7x9LgyzMTVeBwjKXPb+nE0sdgWftCH+q/+4qmoVJtGvsfnSt3vm+A8mrbwlkuyGh0a0PJRqYqAgg9sv+H7DE9NasqP/DlvmTsjRzyIBHSj/F6nrhfLzrpHt091Hh26tjhKN1BrvExkPTboetFArr225GOD6EJ9A59+9jmiGnfAXzhKOPhSyc6tuSm5MlqsNliGFmXqHRUkvVoG4mCt0SeI506Pq+VTDpRENzneE4m0dLKJNuY+PIgSnmXRViMzXds69a5f3x/GvecaMCBn0ULTteCeSkSWKpRvaA0/tV6zloFTlzoHPHwM1XnTyVCOhnZc6Kyp60rJUHR6jUszdEshy3XnHk2uBZPjeh6tZ+y4gLh2PK9kv3U0zQs74o8T033SdI51koT8DgWNc89+KHreE2nnWzA7ub69ZkrDo/H2+qxzvKCNnnJtZoRzkjoEhz6WOJ0fUvENLR3wmXjnpeZ6OsYIsy0cKzrT5KWu4cWPfOSAnvswukbsF6fOnTh4lGccRZP2oR/PQ7WRa26uu6VvcZpafufHpFM269A+aEUPtPWbKMW/3BeN9ZGILnSC5lKWnkfONXL7jZGqPS9xv3HtPjk+5wcPD9YbrOswC15wQzVHz2PWHvo1H8tnpUMgvbS61pfjx1pwLZ+Jf6xn15gwyqNu3FLAaGO/N2zrcyBv2hz4QC8F+hlHqTSWxowp3UCfDnFnmwJ00mud88cvYr7H2I2NXy6kAe3HtrZ3X/XN/9W37n7zt30b5xgCDNRT/EVl/rzqGshl/KoLOcs3a2DWwKyBWQOzBmYNzBp4GTUQW4ebdqyZM56xOjt+97ve+Wu3Xnzhg1i0n9jg0ZU4ghYb5974m7yJbwPgQXx5Y++NuzCaZyYNiNz802e/h8m2dkiY91jHmzq3bCRA5dVX+MuQsL1hxdNvL9OYOTjkMTeixQ4Pj6C1Mig1rDSkmq65ODRK5LedBJZNMfKBOTg6isEtrI9wtkFkf/NQvA0DSrYx1pWNdjK2McebBl6dYr4iVALrSiUt4TyQDPiVfOKsvnJCALCELfiqN5z9xYeli3isy6vjmiYQNi9Tjy2a1de6WAKNQsM0H93f7dan+Lpse+tsOrbLnQvXyVUVlxb6aDzRVnTWUCtddMtlXNbbEJ3CpN2+gc+8dWUuTQ/LzbvjaxzcYdwHhrZPP/vZxXocZCt8cUa4pnBOLBP4QLDELYwOW9uWCZjwZJt9JvLQHfXp/LRuQIovo3jeYG1bv4BXPOB0rIfr2PW6jbG/zxss46DGsdF7M4m3ZC2Z+rwRjWnaN61f1lV0BC5pRq5LYy+3i2s6xnqnpaycmabmscvWdZTFiURj07O/U7d13u1Ns+soJ+ObRuf2T8uNx9z27u9yHi0c86ZTqeFck5eTY9SHeTt1pmvR9qbXzlRxOMbDa1SP73bzPI43eJv229d8Wp6mJZ3Bk30N233mPd/hWXeU61b+gbdstWFq3MXviKZZfTWm4cWjg06Ha5zc6NF16DXdHz98OYEOuP7OEFfRhOgDyuL1kFcPcXk4Rkea5YwbcyNs8VVjNnBGbnqO6bQcyf7G2/A1pngRrPVmufssm6z3If2GHXPqd4ccI+Ma/tCNR9ln7to/8U/+ruUaLyzz5ytNA3W38kqTepZ31sCsgVkDswZmDcwamDXwxdeAt/5aHYtP/PqvLb7pP/uzn1hbP/0QcU1PYlydcnO+xa/4m7n951WBmAcxuvqmvnPZ6kgcb9/b0DhJtEkZGXVTvzIA2iBxrGM0HLEGZCbRB20kaPh12ccn+zA66wSD3l/qPfh1nX2fjnCIHbOJ+FEMJqPGjDYxqsxf4ENDgiRp6hSQD42PLSMB4iQrYyk8DRjlsZ5xMCi89RhQ5M2j/WXQDENKBxnOuRE4IDxBOxtruzv7ccSJR73Rqhkfw041DFXQwnj4a+MZ8CRpFJ2VsWlHt7W+ul6jSvcVzSHdahUWdNRjwpK3kVvt9slHPsegy3i73nxa9xCXybIRSnmsSloYldW+wvuSqDK6jEBpvRt9ob504lTU0gp309fBlKgVYDpBGYITfgZt+1tPyaXF+Ioi0aBHD+pfz4RGuXoZ8ji2+81dk8p+bgQM+bOfeb7OE+qRmfUZXchWKVQUIOFxX4zrM6ORiEQUxqgZGoErOQVzbnx0UkcPleBY6lrx4MaInda5TqH1Dfze8kM5OpTueGwrPAw8AFEtJ4XreYd9xnwJxQEbvB+hR8JHgzc6HvK33sTb533PQfNQoOXYUYUGJhmXGj0oeuYIfXsORGaVg/yKFxEZROLMhQcGj0P8WQf0mRstJXx4AjbOMNp6HvUs6VAJr4yJjtUFhxSbHsXIaS6MPo/yeyRaJ9clOUpklDxf0kXmg/lp/lZ6kAo4h5Pecq9jeboMZ93UuXgbJu0J/XONCMeBfPY3jOeAB1PPWvScrrnd1FmWMYO+oxGw5aC6xJGyH8ioq6gdQMK6VitysOTiKghC4GRH+VUadKuXfdO4prK8Mt/9Q0XwANFruHkwdz4iw1LHyqq+x7nZa8EzUH7QoYeRwjrGVod1r/nMv0fWqvxzvUUtfT5b7+8QZn3SP8bBp2M7JQoMfWftjagxdW+9+TFqUkd3zdBwnHPuOSdGnVbkaTkxHef4Th2F3eu4IyE74hDcvLhy+aPONWKer9/87E1UhBOc/UKFa903zjm/+hrwLGITpXIAACAASURBVJnTrIFZA7MGZg3MGpg1MGtg1sAXrgHv/MuDtXa6+OAvfOCZ3/yNX/spfBnv48b95sYGOxJhmVDmPp0HtjDG+uZcY2B6yEobEm2wZYNkbv6ncJaF8xDO3LYeL/5p3fau29cGkG0dvWWuk8KIsZSp6xAjZCt1cfTjN9ITxtSGTUeDGT1mufuEk46ON8cZoWBdo8XcNnlqmra1TG4aTdLJWMSwFcG/hYF1trO7dfeRRx65xfh72mscbSFh4KyMLfF5dOpy58L20bDmtl1O3W97w4ha2K5P+y6Ptz7F22PMk3TeTNJlvuy6PL7bun2Ja8BOaVjuQ4O5k2O7PTlzYrI8TU3DOWv4af+0fVpuWNeP7abGbT6N0inYBW+xPIiDSpoawAheYxzPesFbUqSHcbyEa9zAY6lLKIcOrESWDfriy4HOmz8fo2y+pMmaqvHA+qhw0tBJdCEO1nGfb47BlM8m+9s7tb8a3Md5gIsI2YeDcvDYtApxzW3ruNvEGQcJtCzb3zDWLyb7pDMcG+Sfj4Z4WvbGs7HuCwdWvNgvHZ1anVwVPa5z+yybxOuYnmvbLDfvPeZyfdou/HR849V5W9NStGyf0m0cnbeM5j4Car7SW53nqvGlfWJeyVK1ksGN7dNX3r/grP76lIapebDc8thjfx/2Nbxl07QeHAxqXObi6rqwaqIdz6mPeRDGeuOblh3Das/ROMMjp5WP1Tf+aZ8Otpaj8ymcZc8FU5fNjRaWlmNMWU8ovaLHeOR+u6L0+lHj4HQEYz0ujinYbksnH8K1nE3Hvm6z3LzZLPyIgr6xs737xPb29rXt7T0R+QRqMeqgOb1iNDCJS37FyDwLOmtg1sCsgVkDswZmDcwaeDk0wM30COXQrji8++Lb3/729/+73/CVX8Ev0/8MdsBjOgCO2L2bm3ItKzbrL6PT3MObeHNMwhgPOqVMGtt0pU+jwrrWUI3x1/ZyVGlANx7HeXefX98bL+ik4RvsjEI6x1Fh3cgS8baBr2FhORE7lN27xjYfLxO/RnIZGcMYod/6NjiE3d7dBhb8qEOe2AQ5ji8f24x84BI3qOIgM9LB8cdEqbkHTssg79LCVYc1pa428Omdb25v+PZLNpJebHzS441f/uYTHJCPg+PLadwXsRpSJvhGxGGIDp2RJdluMpdmp6Zvvds7vwzb9cbVOCovnHHKgL/xqkvhjXCybHv6jEpiYOOMY0YW0VW3ibd5sWxyXRWOWjcJHakukIF/RMaEhjITGaEhnZdBjLVmnxEt+A7ic5KeESGCE/AYPhvlEg8NLYt9bZzHdQHPoSFvY50ZwWfUCB2RE5LUWc3ogcbSQWDWeDvptmB5vBeoRKqs88ZHHcXZI0jGOgURlYmTK2/6o8mziQ4JqTgtYn1ZJMe7vpwDCMkDjuHpvAgVWenmH7UpSwYHlzgzL0b7jMc9T46OQ4MzYrGHDHt77J925qPJhVt90RC9tUNQOqELS7KpE8G/nOf06UAwWddZnSgj5HB9y19FLDKWLuucZUAqb/FqG0sAuoUnkZS0lW9UuMLT+ORF57m6AWtwSl88Js/J6GPkcTjaD+fCRyfQrlw+Q5y8rh9CNq6GMe+j+zqXpuWGtZwDPPLi9bJSyeESMwnfuXpXB+uuPdZ1udcGjHIM/C66kpu+zKuaBGEEHo+DD3rRjjSGXsRxIbFWhKmruNM+zvul/Ky90CjZ9MSKQd3Le8OLt36UKFK2h5aRdIzPdYJxHRkms1lDAw9nTcEv6TaXyg00IkT3WTNVll70Te705RwBMFFv8Fb8lbwtd61DnWAl8dp5XZc2OTeMeEvEGLrzfHe8620L5Nt8R2yNa1hxtlof1uMM5frvdTQpYz0XB9/jPCieWAtcI9QB37ABl3dp5cya6JbzD5QuCtb74nz/8OT4DfvXr72e8m+gGL+sMp4PgEQ46C/XW3fP+VXSQM/yVZJplmXWwKyBWQOzBmYNzBqYNfD/hgbG3XT2ImOH8bWzn33vTz+5fnb6Ye7rn+7X1mPkxnEjg22QNrMaGm0UmdsfI2XcqFs2NZx5l6d9jc9cPBrnpoa13EbWlF5Hb5lr0DjOMf32tB7T7eJpo0RHmMnIMds8dACYCsfY7H8Y7f0opXDi82hehOfQ6sXxtXFE5RRdYM2c7+grwGD6FG8BfMfO1vb/8ZrHn3jr7u7uzwL/SXAdiW/Q9PEZmktH09z+hjO3b4xZttvWMD02QJOxPabzy3Ddbm5qfF1WZlMZb6Wn5qVhAsBH83OZ36bZ/Q3PDKfYNO2frifbgwuvgX2msYCXfDatpsEMBM6P7muc07bG1zCd285yXCbbPXree30JI0vsG764fe9++jc2l/Na4wHQYVXGMNkwktMJaPMcRFrSOF5N2WR/yJsGP+AhHjiKxeOKydQzTxN9Cj/OzcbBYitDnj514rj93S0eNeaMp611gEsjzouWVTiTeWghfJe7z/6pnrpfHJ26zXoegyxxC2eprkHTZqXxt/6n9Qbutq4vx034bvnUY6RZPrpXfF/GMa0L7/jGa5/HEmd6Ll4r+3zpfIAk6/Xo+MbTOBsuuCFsuymOG7xqPpxtudsbvvPgbOfP8MJNcfe4bhO+57lxVF/XSnbhTOGL8rSex5J15w0YHV/i9NrRdHTa1qOvhTfOUIqtiylfXpObTtPsfvE27s51lCV6GHq2cRWBrrotntMGfR2L4rFu6vHy5feJ9cAOnfuYqnv0EbGVjfmbJ/PGo4zWfYzSXHk6ilKYmreL8yycvExT40wfHTWW0fVDVXDzuOU16m8kovnL93d29zPedYwaOUrYNM4fV10Ds4Psqs/wLN+sgVkDswZmDcwamDXwJdZAfpLGilgsPvbhX1p8+7d+y9PsifSrZ2cnzxvtQMJ5hi1dZYIvRlQBddva6PMm/rJR4WCNBo0kj4Yxd2xFGVSunRLYiSFlfwwe9pixX/yBcc8ZN2c2gosNmj3ch2ZlaBPpgJdPOh6Xk74LtstPNIeOQH/x9zDK6+TkaPnYZNEqJ0nz5lvN2nDSEacxpWp8myXRBfgdjnGOLc62t3gzII807W1vPUnrj6ydnX7nG17zmu9+8xvf+KNbu5sfQYIX0QHIyhgbeoRd+DWCQBuHqVnHYWF6kCzqcDofUxj7epy5cJfTZYPUftvCA+XGJy7LjfNyHgNPI4/jcjRM4xK34y7jqv7VmtLAji2L7E3TXP49siatux/SSMGh3oz20HHAgRiJbDH20SgukfZaVRNGvdgWfpw/V2jy1ZoRjz2qrg1sSbo5t0m6Pnp7yDowykkfjyNcK64Tn2Q7Z00lpVxeoDjHKLYe0886SIhJwkyQYzj3sv+QZeRAAtY4iNSz81uCQNDIH2SRuPNgYcxZ5l3BoKdul+vARTrWhKM15B95+NpiRx+euI3YpF0ZPaaOCs9lnRp9XvvGTKPFHFeH46A3DuXLWiNn2IWUucOwP2VPtmPPd3i1Td7Sp2QDr0pwHnpeGlH0mYoKqbWU6og0KzzgA6f0W25hxB2njgsFuoFJRM9KdiPWPHB9MILySH3+BIfCTpI0bZE3z2OnwGR7ioFXRrQ4GZv+lldHDolrcdZnHGL64VE+P1soKXhLP8Ixu5CqteF8WZbrxl954RTe9encmWetDj66PWtGfuWH9dBytr59ktx9x2p5Xp5ZKehsqvNHUXAfwUsdU+h1deuCIsmjUWZWXfsu0ZwD0bu6X81LYIEXxjcXH3MN9rFInzWUlu6xXquuLQ/YyVxkfy8G9veLp1XjKz2p9zrkS9mdSriPsqbXZXny8DtEfQurg7wcZeqvrkfiyXLwg6TE0a3nq19ezqhlcg/5CC7nuNDwNVLrhbW3y9y//s7te2+4feuFXRaulBkXZkqZA4+Nc7q6GqjVdHXlmyWbNTBrYNbArIFZA7MGZg18qTXgHXm8Df5K/r6f/qnPfvLpJz+0tbH+Ye7j7xABxRNH5+vc8PMEGuYNN/8amJePvpmvG/4VjMLYNz28h9f4sK0NYZ0Kpsar86nHTNtta8eUsOIqo0saOCmUhqThdzk51hSjw4gAogF0DGjoemhUykfTbR6yEfuQYfB3zt5khnsdMwYfyakPg2EqnuETW9tDd1sctzbOTz+wOD34ew/tr/3gzWeffts73/ZDv/T93/vdH9lcP3+GcXcxhnyeMrTBFd1K2zTNu9zt1j0ce7nPtoYz77ryTWGtt+4bRnjbum7+oHLjaR6mdLpv2qZep2mKs9sdNx07bbfcY3QomNrwX/Iw5C64MjTx6uLMYma0Li9ZEfZN6Tmu9aFh7dHG/RROR4frIbAaxHgJXEO+NAI/7eIej+eqW51WOk3dj06HQ9oskIJv0E87ZQRMn86HOCBcBx4azPYxL82HvKbsGhjwS7wUooOKJsG1Db6hf9vTp/Yo91yfx0l7snjoOoEo6De6GQ4L8fb+XvIqXcea9yHMNC3xyv80SZO21rPjdWA0TkEbp86oooOrIyoY+lnKMPQ4xjSZ5q1x6dgqvlv2oR8AprDCW/cwyYdpuna7LR18NK9d77zx2t+y2me98U9p9bjOe0zWxhhnX6/LXKOKzQwpXIVbB0voo1mT54ttxXutocZvf/NTsA1XvEp/NQ+Nf7VuxHMhoeuW2cuvjiqTG+F7xgp/mfaUvrDLOrim9abV46XjoYPLNnntvmWe0wYnGIx0W4/pcdIr3xQwqMx+k/D2Of8e6tCIVOl4NJwwXRaOrjjHlt8rXPritGT27HMsX045UtSJRV08attkeZqLn7Y1eIJwbS1wfHqyS/sb+B56A527wjccxcnqsGdOV1kD8x5kV3l2Z9lmDcwamDUwa2DWwKyBl1UDfdc87JZxG40lYIPBTOw9dHJw5/avfPiDH/7yN775H1vb2vwqbrqva5Dxy7UOMm/w142a8kbfwzb3GdJQXxohibSoG3YNhfrVW8dCGTLe/2OOxBBwPC6qlOkmWdahAoRROOIt/x0tZTTlDZWMq6SRpBGo8dJGXO1B1nVp1IHDAn7cG8ZHKzcTnWV0jG0afvBoZJpRaWzOb9spPOgoOzZKZ8h4enrC4y7UQXtyeHS2QYhS9gHCKnQvKaIYDnG1ve91r3/879+99dy7/9p3fOuTNz/zqfvR88bm6f0/+x8fPvTq1xziH0uMiPyb1J80IBxHwiaaCd86VmjTUTBN9sljpy7rxEkZ+Db0uq9hHdvy2DbFFZpL/YJrRHMJ13gyXjtM3Y7+NvCEMzXtnp/p2C6bT/fqiYgdVUOl9OHCULcVUVKRjcYsrdaQ9HpvKfUUeZQ/SrdX3TrHyD1k6/281BeSMSYL0ArQaZlYmtCnlbMA5K51HEmsG/nbIFrQHN/Y4uiQc2OTPe22t1TNWJvgg0ZHKaYjVDh/6NA0ll8jjVz/YcO6enB+xyFk5gYBa9rHOGT0T12qA88tI8DiFASP59P5Ou2iB8Z994hqZI3hsDDCTWSUH33oxmIP3tfWDoofuXE9uq6BMTpHhdRWSWgjrEETOA/1Kpzt8uM8WTcpTnLwqTvl0FmmAwagrJUVkIjrbB/DQMC1QPn5s5T5zQkBRCMHV9ZcBnmtGLSBl5ay9Bz3kF570T8KcoTXs8hNufQddmQ/56A8mIqHlYw6WMTHi2lzPWTTxiVc4J1rZD0F0Dx+EieJuQr9QIuj12HJCTcQKzEdZ3RS6bXWtHMnv7yFOJypJ//amTzQJjovdJnAXlfqpVO/5REOwMV12z540Qlc9EqfIM4QuSy+S786nfyR4oSr2jFrxrmYOqdcSmKQ13xnIEunmht5Bjd4cioM/NLRyRR2MmasRZ1ooHBMrjFUzV058isN+4y8kxfPjNDxqjuu56Lz8Xn9iUZ8mcKn3xGc38qfSGD25+vzwGXn2oZc5kX81reJGFZ+nWkmpxay1NHP4DNz5SxJin73vRSP52ZdC4Iy56gvnpFfleGbcoh25muWd/7atljsEln42oPDe69F6J3gy/cuTjQvVArmtWpOV14Ds4Psyk/xLOCsgVkDswZmDcwamDXwcmgghtG4X24Db9CxVZsOE5oQmNP123u7O7/MI4Jfwy//X3eyvva6Qw0Ie0gaGt60t1Fih+W0c1Ne5XL4+Iu6ziWT9IXpVDg0BjRbanx4BK7HCJvNlr3RH9E3MXTAE8Mnj+AULceabI8hQ5byaEsEwDD0dJJtbeN+Ii+HWfFW/EEfB6CPbB4ckWvscYAfP188We4V5vvgNk7OT9mPvOjizXvh/PTwMxhJzz3+2MNP3r936yd+8p3/4P/88bf98KcOXvwMXJxq1cD47s6LL3x2/VWveQM2GR4VUvPeuW3qp/WVjZltJJXcgyZ1xwhnfrkvAy59TGFaP4JcxiP9bosjY+jX9lKDczMMc/qEnRpkTafl6Lq0HKeD0jb7u6/lEKZTaOBDEcayqXEu4eNQvShDAF3UjMMVlKo4TK2rxhfe01N0dB4UbqbMpecKlT74goNy60ZeNIC1uX1K8oBN79fXdwqbVq9rWyT86xgBQZwnAoireHH+pEKbSwycyzScKWwESJ8QpGSFW3x5xq3bM081H4HAMj/DuVQ4pVPOZ5y8MCwuxksPI/+h/f3Fjs8fDzqlL3BBMHxKg9R8F+8tg3nNJYXAoOklrON0XdRLAwpWx7mt0Y94+dO6L7r2yBq8DYeR0YA+0ipd08rZteIhHZyTuW7oqMCJIr5eM+kfH3ZHR4Vu2vWSsjzq4AxvwF/GmTqbu4eOMnlOTrDYr35MkYm8+4OTeueKV+Vab4noo7Ee59ZZolz1aKP4oo+hI8vOFwBpd/WzQARLCl7HPyDZ13OaMs7+bhN8pffiK1QY4zzoGBLWH0E8TZVf55hphaPqXj/8bqhzrLQgjHM2pdFjzyPbCk5H7QU+kTm45IHVNHX6hTbtgbdX5uQZdHGMQcT5aHz1fVDrxcdH/RFli+8Nx+kwq7lrPkse25Zz6jVngs8XVsiDM6B85zjhkitv5FDKuoa0HmEm9MTTuoM/k+0oNm64TX6ZedXv/r3/9Kv/2X/x6/Z+9t3/V8mgl1ME6MFPyMzpimtgdpBd8QmexZs1MGtg1sCsgVkDswZePg14w58b5r5prjyf3HwbGKI1evj0008+y6/pH8WQeRKj8HdtYtidYANwWx4LL2+rnNzEa23klhzkRh4YZuGN/Qn7CpmLdgMjw31bNI680Y9xi8GgEXBIlJZwbViUGeltPgZBjNwyuk5Pj2JYEUpUxoXGzkihgzEcw0vjYBjJZ/DA5vjLqAsNlt3dncUmxo5j3N9na8s39/lmTVxWRI7dOzxa3CeKzGihQ3L54LG6dYx7vAqLUyXBSllsw8d5Iu/OXlzfOH/f6177+p88Orz9oe/6zr/6Wx/5uZ95BqfDMxtb3r5qpA5mcapd393bZ+z+EQo51nkxjHiNWWlFbsB1FphUoW2d5Nu6ecqXDVlVXoN6SORzjDo2Oc55FTQGN3njNGJBh0BHZAmvfhxr3rysD7riMhlF0eU08CF8eBz8hy7Gsbl7gxlB0Z4CnZiCaUBmLTQS9BPph6ErTpNzLR6pN++Oawde6VPvmtAsYLBolJbBzRi7wvtwOqgP6msa8NFTyaXDTMN/S34DX9GQRpDJi/R84+F9fMHtFAiPni7igaYprgvnWmmUNXk0LSM0gX/oybrrwrnotGaEis5a/sKHMA3PjFUCT5SoXpSn5qskKfmMpFv4FkvXnkrAIaYT4GHeYMm7OMFOpGXrdsyf0xSVQKR1HRb5kBfnwnXU0YbCVDwTAwRMVrAVPSRfNVea++4JFbyypt6UYVxHRqwO7ntOv1wP1EnhiqzBXh81P4xXy+CIcxA9mHruLGccaOJMiRrRqR0kr1XCSiq846Cp6MO6Fji3rrPGVxFDaBtVej2Z8hQegK+2Ohdci9ZrvzPP95Yl5JcfRibRQx0Y+Ok3J7qcSkVjHeTHA+FgwBHRIR/h3zVUdNfXtoI785/S0InrLGmsHeSNbEa8wasRYcrrOp7Kph66XjnzyDXU8yG+YJhUgpVj0euHNFhywKgH6bhOMl5+Sa3XqiErY8TT8K4X580107Cuc89v68KKr/VQc1fnh/2J/kIevw+3yHOuhk+i8+DNiDnlrYiyYmo53/KvE9nEeSQ+5ZOe8+g1wTZlFKqdxn5fCCctz/HAo9/it3LxOeYMx2L0DU/Fm3hKHtqzRZvjcJjuvvZ1b7j+t/6n79v9u9//txd/8c/95wKWAmFb+YNw6JXanK6gBmYH2RWc1FmkWQOzBmYNzBqYNTBr4OXXgDfU3ieTPTDpOIjFgB309JO/uTg+vPfU1sbeL51unH8Nv6q/+fTkeEsUuVEXWe7ZMYiGoSPS0BgELGMLxECwz+gHHzPxhp3NVAK7gZHuYznlYBjGA+OMmDBp0oRem9r06Zwzysb2NtCMLJEeTipk1OHUhmrtH+MjSUYCOMYIAY15k0aIxpD0dY6J+4iosUQDYW4dHh86BhbP9NNtYZRta4vyZKSPmT13fHz/WR79+dTDD9349VsvPve+v/O/fs97fu79P/XRu88/A3IMZYyp06PjPbmBXIWLUdjd3tlFwn1w4YeB95JXzcjWSo+0R9WdS1s5h7zRDfU2otpB1e0ZCz7rnaZtrT/bpjANa277FN8UrtsbLs6uyWDxtxPL5qa3LCOHSXmqL9UlTYStBj6bVufVUf0tUwOLzxS50GnryyXuqpJWtzVc5+IvM9WWMRdVXOpZGNdoYHES4i/Vx7S4f1Qb9rshXR4HDf/oHnrB6Qw7d04H8KCgazipuo32MmxpUDyA5FXnU6LLwot9Y4BCWU7VwcBxjMew4I015Bj9ESb6dFIEL87bM5zBNOIkXl+86pEbrGvOTR3WDFBPOnHUprIK17qjciF5DgnzoP7L8+NA4fByhFdYinNjGvkjjCR1guCuCG7xZ95GhFvxVLxZjtzmjlXP0hhp2SexkeShcUx5bNiGi+QDtnloeksY6EYmGhqvufwK69HtspA+2kxT2tZ7nHOlk645bjivYeX4q/O2HF4lqyL7aHnSciDXuUG/rn3d0fM65a36omenKHKXQ8u2Ti1T6aFk0HFlcsWc8xKNnk9Xv/y6Gb+p5VAyy2MYNeaXujTl0xdS6AgUb42p741+dFKJbRc+eD3L1GmxASOOr3rzbj8zQrty6sTVGVyP2NsuXF+zLAvvjyqm4BD/JNlvk2O4ioWfdkDaJ386zngwEn83ZfKxQpEbvodsBVvnkN9XntZxvOGxK9mXRM/5Lj3fxFmunilfA+Hev/B1X8crmXk8+vQYcH/HmdMrRQOzg+yVMtOznLMGZg3MGpg1MGtg1sAXTQN9S69d/HlSWRkYG+986z9gX6WdF7/hG//UBx5+9PE3c/P/yMbJ2au5ocdbxIb0WABtlGgYuG9XGwMaEXGGgScOMfcV1giKoaCxUrC+tQ6IsONjX7XH1zCUh8GDRaLJAQy5QoiTLI81xvgAnQYQ/i4fywQcOtgJGjwYNb55TUNCeN8qqdEc4xI88pkIhNPSjpFjPhF0zHFwfJRH5bBddJ6dnxwdKzMGC8SV5ezkMycnx+964vHH3vXiC8/88vf9j3/zM7/w3ve8gGfhs+tbAuGN0MuW9BKtE5yzsbe5sb23vn6Ad67h9Bu2wa5RpWFUBpeRRNKHcmQwSkO9L3Wq0CT7k4+65Z4XYYOjYc3Ry3QvIGFM8iGsY1c8lRHYjpCGC/4xRmPeusk8fcFZeK1n3TAv6WM2q63kZVTmL5I4rlAhFQ6bxj3apKHhHD6H3NXm/BTtdgrEUNYYTaSHxm4ZnVPnQ0xgcOuw4s0JIV1msVgZMeRKRbrgQqOJlDFo0rXyws3bi3sHR4uzvcKv4zNOyziCoN+OC/GhX+lk8RrFZULIzCmghon0uZJ5YU461TyhkFKKzFGu/tIrVVGrX3jsdVEhUbWufB50bYOIIoWEv32iKq/vb8NvPUp2xvkkrjjmPOsS/WKkXJ2LoSN9UuvGvMvyuI4D3PmWs8Cz1h1iZKb96jrwObkBQmbbG4djXec0ZIbz5kbGmrfzq9dn6URuQDPBM22/XG46jrHs0fhskx914/mnOitSLIXwEweHqrff8YAGR3QvHyJRevgdcpnzX+uWPPQKMGVHNB+Oc524dJNGoZxj6YV4/uluHsMpuEqP4nKtxkkDrvoBoWSVl9Af6GUXdHDMtYXxS11AP+eZiwqARCKP9dhyWTXSzOuD3wf+8KHqVErkgb9Eb0KTsz/4lvjRX5y2ID+h36irI65xyuSlVH3xtUPdVLl07c8eXmPu0s2H9DyWTuxBL3zAKJcf1lVHevHYpE5YnWDgdCqc100jf8PLWBPgPRWnayvnAnhQh06sRJ0NuuoJcZgz13+t5/DquEE71x3EyPUBZ9j6WP/qXZ3Ig8gzDn2KJwn9Z19O3vJi3X5+4NkH796nf+tTi/3r1xf3br1QsAEoXSzP/1XPXLpCGpgdZFdoMmdRZg3MGpg1MGtg1sCsgS+NBjAXipD2TQyLB9Id3hg8RhgLP/ven37xP/j3//T7jo8Pv2x9Y+f3sGfUq48O7mt4uIP3BjfyOzFeQSVOb+wbt7nGiFa6uUaTadnPo1Jhw0e8SG3QGsUlvG/+E58GtDS0H9pgs549aJBJqcR5xGOQ9UicuHAmxabGGebm6eDLL/rJY3lAAzNR5xPOO3ZVCy2dYweHx4v7HIdEkWFa4DvK40IEqK1v8rgTA9Y+uX52/PHt9cWHbx/ees+P/sg7fvJHf/RHPnV0+ybOBhDgdMCx4HNMejzwtYGgIsdktRKej93d/U3k4742my5HBp2K7byD1SRlUQ8wPAaXvOqgddw6VW/dJrDlaX2JYPQ1vDRMDSu9y232C2+f+YOS7W3IiWuaxNf4Mxejc9re/dNxtsle8eraaKO2eHD8VD9L3qY8Yux2tAjzu3XF2gAAIABJREFUUejLe5SyxiqIBw3pVbSWnZflaB7N82ICdcVcRHbG3blzj3V1cdwShzppOkPHrkHWgKQclKx1kjo4Qwt4U+mh4EYD45wTHQUUB0yV6lzQSxFnkjoJPVdduRkijzR4dHmP/cf22IjcRwRDE1zpZ1w/cmjeyT5T5637HmNfO1NtC9zIe4wwJqejx1dLfXZb47TuoTrMdfyYel02fI2u9qbbl8CGbz1Px2QtAdD0hM1SiacnHTah0nF9q2WYtoyBiLl/U7zhAahu63xKTyS2T2nTUvjGlOfHgFDrj6JzWf7GIb7GiSQZ1I/AWrEveqjlFT2O4pKPHi+NXO85n4yGkrf2a1akWCmD3uARxGu2By7n0PYjOHB2iU/a5rUXl/Na3yPC2T5YzjpynD+q1Jhaozq1gg/8Latj8+MI4nqtyQoZ55FjW4aWnSspY8vFYL+Hmoq8lMMHSDYQ9iwOStv4vmHt+Yi4V3plHmdx6Ts4Sx81FwB5HULfncrxOdrwd+nUj4tT+qyhxuqPPOqyvkO5BhKynEeQpcE4+OO03b7B97Pfyf6SoLJrsi0EV1Od86uogdlBdhVndZZp1sCsgVkDswZmDcwa+AI10LfnK0PkAsJ4AbhHj2Hj3fOD4LUCbT/lfut8/cVPP334U+/+yaf/4B/+Nz6Ip+djOJW+mh+72TPrjKdgCtHxcT2G1Tf+MS64IT/OfTro+CndG/R2kLVRYoSBZlN+ZR8GgX2HOKdiCPk2NsZt8kY9YbFa4AsDgoiXGGPYAMK5/5c9GxvbC4yEPBomD0aN6WxqehpSGk0xO/gwegDLQg7gzb1ceFMldO7cv0fkGJFk1Nlz7AxHna8ES3DBxtrGx8+Ojn9gc+3s7T/0gz/wzE+/68duLs6PPxvbSn4x+samzyGjgTNSMT9p0KXSj4XKg7LKa9k2ijsMR43E0Z8ScCYNUw3d6GLYXBqZGlji6iQeU2Yr+KtPWibjEHSerPH4aY8LH+m9+GF/z69GY5eTo1n7xW7d/pKn5WqeKo9mYmg3Dfmxb0SWDXDfXGezVff4mvIgful0sq9pbvj4EX1uAr/iR2NyKAuEwqKu5HBbPNsuLY44QQbyaBH82WOLtiyI0aezNiuLMJJbd24TCYkemJvg1zHMOCp16DAA3situE5regKrjGrQvzAh/nG+srjiiMv6SDfznH5wOceeuuHaRmjH4C6HtfIkSjF80Ov8+OZKuWajfg9OnMW13b3sO2ZwCo9Tg0Ud1gs2ej77fBblUteeS8xlzUXNQTlMAIKtWhfKHY5LPruoexmpPZq8HhTO8DtcDvSWbHr0THFQDDjWhjq0J7rO+bZy4AW8kMKbjNhSdJv3znstF8Tqs3hEpjGf1h3DVSNARrKZij55r30gbKuoKPsLrvWicyXXxCGXDvvWh/gsm3z8TwHlr1PgmCPP3XTy2Y7ptLjWRnJu44hhfPPoHPoIpnjEIanep83orawLf7iAt76eSF0ePB99JD3OYWDPexN++p1/hysX107WEJGIvAglOuA0zQyP89Vrv3O/4blCrl5c24lENoqKP/HUDydcIcHrDwjqUTruZZl5QFbl2OTaIH8lY12nlvLCG5eD9ItT9Zzp3AIeSRgPAEnfr/4ljx7bkahsPynH4dfvnUQwc82vwTU3Rpdt+x0Dwp4tRGL6aHP90Y/E6XeccEiBTr168Mdk5ApuH99rzhOfGafeaYa3rA2FzqnhdxzfIzvo5NG7d+8+fHD37vOMyDCHklwMQ8LU548rqIHZQXYFJ3UWadbArIFZA7MGZg3MGvgSaUBL47e7XfZVeb5uD6Pj7/+9/23x+/+Vf/Wj52ubb8PSegjj4GvhdD+RVdyvY2R4M+6jgXkE0Zt+H3X00RZM7whlWyfLGikaOWXsWD6JsYKJEqNB44THF4dzjL61Dfxodc+/iQFi0tBITtgW3Tw+uZ06v6Kv+XZETC7sQszGkTT2LLqnjdaW9LUxFJM3dcYhdvf+IVsvsbsYcWO8CGyTx8O28qa/87P721tbv8reTD90897Nv/Od3/XfffSTH/8I9HQinGycn5xJHMbcWtldxD1WjpswdvHjHD3qeXCzGMuRF/bUWJS10hltw96V53aqia5hzB2b8RhiXRbGMeKPASYcfw1vv7D6jBJhRN2+ppe+zFPhFl58tmtcmsxtc4ztcm/d9qZju2XTNBfclHHkhWsF13Qaz3RsBl76uIin9N98Oh+uN2lqjDffQcHacMk7XpaaTteF6bZp2TY1ahJWP9Gt23cTmbikS/tyrDpzHdumjpwX9dIwtFkOvqG/ZRnH0BIPjT1fDX+hT5wDl+0a4OvuWcV5J33HalifeJ669uIgO1tcv7a32N72zaIsTcYZ3aZc4jA3vYQObVkTGPfCtF57TOcZPGAt2164KrrUcc68bZYHOUGrDRm63LwUvRo/piGw3S+8ZWdpuiaX7dAK78D0mMv14tERU54HXsabemxo0WYuHlPLY95wtjc/Oo2KRuer9ZSxkEh/NS9xZL/IIbT9WU/orfFKo3UaujowgdtYrzfHii7tJcLgWR7sqbnHDTR4K9jasF7MDiqGer6l6xOR/rBw5F6TXIfiUKJdp3JFShYe+e03qXL5rX6vyyTrOsciU5rUI7RYi7UuiC727bfI49o12a4jr/qLRrcXLfrG9dh1b5so682UXq7BEefYar33/Nmnk0yfUz6hpVPPx/UzxVw71IsOQZ3eOsd1xnmtCW3HS8+EbtEw9eKx1ol1GpTPrxClz1oXFn7cnkDxgVG+oKHMd+ba9uZOvkthfWdrc/0xvlcfA+gWw0oogKWxpJ/R88dV1MDsILuKszrLNGtg1sCsgVkDswZmDbysGhg/YOcmvwiVAWe5bqIv1LFpvAs/X/v1j/zy+X/4p/7Ep//63/yeH97Y3lo/PDt6lK7f4zjcT97ZYxnwU/caLgYiqHCOrWnrcF/OPb/7yRzmBj2PjxC2cHyYTe+56TeCgrdHYuRoTBkdIEkjK+4f3cPWMPLgaHlzr4EvnxunGwRpYYRsbZ0Pe4H2GIbnOLHWtvhp32AxI8+A06bJOKIZEuxxZJQXeLYxahx3cnyWvW6kf8hm5UdH7IuGz25rY1uFYCNy63l+8gEihr73zgvPv/Ut/+23fermZ56iS4NJ81bNeuRXe3Npmn/uhDvx3GfaFgjIB5v4R06MMizHGqqM8skH2MqI2kYHFVVRhrAENAz9exDBNpaDS1jktTxNeVRVGiaMPRF11JVvbezIlOZHnjwajxpQ4hUfhb/7RVvlGlNjy9EXyy881RyJKEuKMU1Do1tDuB2kg9P0t3zSmLY3r1MejBVRvUZllEopu1CGLLhORYM0/pEzD0Z/WNa8rhJl2lZj1Cd11kgZsYvFXda3Dtdd1q9RZqf3sVUlWANZJSBw4VLXYRGdg10N2u4cKVcixRhnBI3O6KUzLZqGN1GKV37F0/M6ZBJj2qF3iixZVmG2NKW0kAJ3XhixODi9u3jVozcWBPwsju8f8nbWmueKNsPVMc4b9SFejfWpfof/umTKbMi3uoQ2Y5TJtMzVbLEfXOkceFMWFpisP3kRPPLiDpCJ+sC54j5qCMJY9wFzntNVYgaH0FlDdmSsLQMfPEpDvsRfNFb9ymhb53XN0UHh+ILjXKZczqTouXGb8yOD8xxRyeXTlPUCM02vNm6v9gAIM2hbF87zEenSjsSMBtfgWfcKl+vVcmq4MU9e/HwEXZw1d/KM3DJmzlP1XMCRayiIdp1aeYwQ7ts55hgPz3chPU987NBLrWN77zGjx5y/k7H/5FK/jJSHrH3Gs9d8dO+bX8sh65tQi7d2CAGW+XPj+oqG09FXEWPyJz/8miFYyhdyZO41J5y0PYQ/TRRlhuV7wNLJWMjCmCKvS3foxevTmXycSI8O9ps853F8I5bX1jjX9bShGx0WkMv5DTQ8cCGzjSE+pqys0sh+ZuGp5MgQ+tSl+ssYEOVcEt49A5lo9eYPUa4vvgi3KD8K7CMQ9fH+cpBJWGZcKnO60hqYHWRXenpn4WYNzBqYNTBrYNbArIGXSwPe83vPXHfMq3vmNgaaLnU6Y4KxgdfZxm98/FcP//Jf/Lbf+qZv/pYf3d7afNXxyekRr7P8Cm72H8Ig2sUE0VTA9se5pKFpmRt4du1anPLIZD+Oc3ZWRqQwvmVLo1WHj4eGpWS59Y8Bd3JUjjQNghh0wBg5AAEMYu/4HVeGE2QyVv7FEWMYOOk41jdTkp/hHJNNfA9r5wc4505PD309JQ69s/PjoxNAeHiIZw3P8cKd4jjDOHoOtn7xkYdv/ODN557539/yl7/tZpxja8fX9f5hwtwDnzg5zEzq7YFponBUdX5yH2Prvqap/JaRjSATI66xKBOsRU+2RU+0abx1shx5R5swtpmbpuUe0+3mGuwAB771J031/SBcU3yW2wQTNuOCrvA1bOBo1zFp6rrl5rPLOoa6bF/z0Ljs6/HTsRnEx4PawheOAmV1zXVq3JnBib4gkLWsbE23aTq+jOJyFNi+tbNYPPf8i+UwA48GrP7jdZ2sGMXScVPu4CrxPGl4/kujmkRf+JaH0d9ydK6hXuWCZUglC4xr/hJhJi1xO8YTzHrAlL3mQFwnOAp8c+CN6/sZH8eee/DRJp6sq0Gm+ejcZstNt+vTNsviMAlnOY8Ds76iC/p1dFDpZRSczldouw5Harw9TpjGaV/3C27ZZL/RTF02b356PCPT70ePM7d/inPVX/NI53Kchear88bV51QD9yj7g58JD6w6oM3xOQBs2MbZemlcTbfrPd66cho11XLYVnRWvFpvB0z3q4/sM8Z6kW6nabnG1fo459p+wj6Qhzxyn2s6A6Sdazvjm36cPqDzJQ36jIy5NcKMKolrNY0lN+uFRn8YcT/KTd6wqpMuv34MfsTpupFOxkz4FFvkHLld07qRbtO68DoL5dfrA6sKvI4BN3zIg6vQrxD8UYtD+DRS7MRnVMdXALPG+TYccnxVGe0LhvAmrbrO92y2/uu8ALD4Ac5zX9l8XJ/LVZxp9iujsiozusgPRbaTeCfN9iPb27uPbm3t4Cxjo1ATpKfrOm3zx5XUwOwgu5LTOgs1a2DWwKyBWQOzBmYNfD4NeHPcN/SfD64N37ppfylk/yrdPS/Fu7ph5+4cV9IJtuz64j1vf+viz9+9/Rt/6S1/439ZrG19/Pbt23/k/tnpP49B8GaMjQ3feHeu0wBD4sh9bzRcyDcxao6NDuPGXqdWjHUtD5JGsjf8OIuIjMC4sA2HgUbRFuNj72CIGL2yYfSUG/HHOMBo5RHMSkYp8MgL+48p8xHRO2cHGjEVcSYSoxuMbODxlzMixfBsaVvEcCF4ZG398OgQ2wgXAXLgxsBQgpO1tecPD++/4/Wve83f/c2P/8pPfPu3/ic3z+7ydrC1YxCeHEIMoMRf4POQhsaQqfVnvcvpyIcyYgLxhMzxAT6gA8Zic/lIUhxRw3+icVyG+eAzRqR0YjTBuwZUISyjSb12Es7k2IZrI9L2ab91YeJQsY9Do0qYZdvANx3XZQ1JBTJ0JZEyjoOuqWFKBvlxXspR1Ht5bbUc6CrGKN7P0NYwBZf49e1QCU4/YjwOOk2rZe26uu+onliZMWTFEz0Ht24padY8sWcdvBilE75pbopGrxnZZRpZPZ6FnEsDNGMXi5u3fcKp9KeDQVeUPBlNGbxEO0U7mS9KyuX5oB7MWYHZlHsZydJrQd1xTg3dgjDRNJmj1s3QSfHp+tHZgOnEOeg5REOE6jURflCuUS27vHXi0Rs3cFgc59FLViUyA6+3QPwqI+xaKJmc88wNdWU28b6LJZ12jtSclN49F6WLyyM6EYdJMsLRm3rNnaTVe7XZwfIBTllqPtpBYl/JA+zQQ+q0B2+xd2GNRg+KKF3Xr2R6nga+4r1wF56seOT1mjZoskrTB93oQTxjnppzr4HhZ7Rn5UDT654p7IXvmm/PD7DTUT8YOJeRGH1Mz2XHitdra8trmzPi+KyZsaa7P/lER3EKAe9bIp0fU848dFzXYdvqUM6ck7aAw6Sjy70ovcY6Xr14bbdfeA+ZrzJOJQb4A4rLXQdZ+sEjaXEbVeWy8FH5bUIadSwVLnAC11GtlnlxCudtrSn10kl9mXp96iDt/qa3gi0enH9ZFa7eYusVQty2cVhD/4ncUjZ+mTk/QvM67pBvyx+AOOI454UtXtd3eBRTev3GTAWbXidd8aa6DpWOXAxxaKdvRPHxfRa9+d2Kd0yHoTrZRjfoh9+rzh/m0daH4d0Isk6FvGtzfmU1MDvIruzUzoLNGpg1MGtg1sCsgVkDn08DbXB8Ppjfvk8za2VICP858MYs0NhZrB1tbmzsbPz8+999+E1/5j/6xL/99V//HA6oWzilPrW3e+1N3KA/gnW1j7mwd3pytLm9vrV5cHzYd/7n7vpykh+8sT6xJbe4sT854fFJrCgcPjyhg5mELwE+sFGAZbd8Hls729naOsVgP3/qqacWu3v759cffuh85/qN84N7J2ungEIf99L2xtbu7tbZ8cn2wenp7g6JSLEdYtPYL3lr9+jocAe8O1DZPjw83NZjoby+REDDS2NIRjVm2H0Ml+DZzc3T06cI+vn53Y3NH3rvT/74W/+H73rL4eK+ex8fXoM9H4vEO7fSYRlcn9cW0dqdJLZIPzlKBBmGXBDJkwl1BFacqzaaRr8wthfNKrcctvXRTpA2ChtX0SjctnlMYYJXFobR2fDTvOkH55Cs+REu7SPvdnN56nrDRf/hw5YaW21V788e3zDWm4+GmfZN27rcfOUMQOsa5LZt4pTT+GznTcObN50umzsmuFSTMlHXIasT4NnPPuczVBkXvWqh65yDmGMiP7wXHsdSsjp0vuxPux0cjDM1L4FJC6jHGh4Ahavp0KjDJk4CLXz4cHlhugdcJ4SP7Z7zUgofCd3fI1qTHvnUXxe+Alm05aYdDpFFkDEPA6zkG5WWt/jVoLej12gB9fxPZZqWxTFNwtc6QhyY1LnTqWDH3NBovfvb4dw8TfHWHJSem7b9F2CGnDrwu898Ci8fPabbl21jzvscaH6cjU41puRV/TrJdAZNcU3LjrOeNoaZi7/SCm/zNDoGvjp/4hxjXNYqAA1r3rgsZ8UAZ7Su9dCFd3xi9KFnHFL+MOKPFfY1ni4boWby0UIdavjFWEvi0alGZVxvfPxQh5cO2+2drVyjHec5dvn8DA3Hkpqnyj2Xq931HhnHMrK9D8c1Tlx2VivhGCx+bSsnd5xwoHRs6KJmX+pidLS60yl2gqd5zf37fBCWsm1HPIq5hQNtmqbrdsq3MOF7nGSInK8Z91urx4fRgdcbeMCZmb02q3zK7wzrD8HHQ4xwkzlRmcSwrKRl/riSGpgdZFdyWmehZg3MGpg1MGtg1sCsgc+vgTZ8JjfyFwaU0YulcaH1cmWYOtzkV88yIqUB+15+OGpsxpDBlYXDixvvn/uZdyx+7j1vv8vP2O/hZ/OPbu7u7/9L//If3PrGP/mnd/auXb92cHR8A4Nkf+94OwE6R0dHpzwux5Y0xJOdnZzhv9InRMAZzzBy+4+rCDtQ/9naCY6eU9p95PBsf2f37OmnfuPsv/kL33J2/zaRW4kYWXe7lcVXftVXr/2Z//K/WLz2y96wfu/ukVFg21hzuzgLfOTzMfh6gt/sH4eX1+CXewIqrwXvazAgXmVkio8CaZi57ximUIww872t9ScPjw4+cG13810//rYfft8PfN/3fGRxxqZSG+j8/BjFnh4xHpVNbY7Wd+u/FXmxvlRrdSuz0WMH2IgEU2AAAYBazjHEfOHB0nnX2EIFukbMSL+jEIS1buRFjOlhD9mu8eXxoCQ9+5TEsklj3T+jaVK/IGealjiXOgA2ZQzR4GNM5zUCvPI3cNonb8rTmrOt2UxfjMBh5MJg8AOcPgA1eB0zTVOaVS49BUbDlb/wYU5jxsOX+zaxRuIMcJ8g0UqnuZvSaYeBON1nr5PtvlUPP9Pi9q27MFxRPkQkgkb3cPEq3vCmT1S92Zx1TZ4y2dCne0ZF7hoaUtaLe4irI/90PNCuU07BskcTQmRDftbKEk95hiVYpBhj9Nkx58I28l/b2Vm8+uGHiTTj3IA/dSxK95fSeadeor+x/iKHeoLfXEOkLV2ZMIV/x6hPOR2Jgm2s1sDnbZs0tJ7VZeQGU6e0KScpkWV0RRfQU4f2qAfhjLCs6CVjQTOg8NEevBKX3liPY2qELD8mOEyRBfnE2Wsy8+c46WbeyAcMUhb+MTZIRlm67v9lsuyRWolU48ArzUSIwrnXJ190YlTXSieQhuHgGBGRy8jGYK+P0qWX37AavNWz+nTvKufYsDkdVi5JV4b0HR9dkmd+xzDbdYDh4ko/2MOL403hn/XiG2SNJJRPHWFkLqE6r1wvVPwppM6zGrfB1lmuhW3Oo01ioHZ2vKRnmQ/cjpe3lQ6dYDUpnd5PjK+YwOuIMzUNfn6JvM63fEaHysp4fqUJbNqCP4/kp80FZiRl9n9jnGMZlHm3LH6dd/EUhmDvJ+kMc+7HOYY+xnpDNaFduqrxwQMN6bswzCqBlzqfCprkdR54tgYgYo952GAPNBxxnKrr1znFrwNkuB0Zh+JVqYdbndMV1MDsILuCkzqLNGtg1sCsgVkDswZmDfz2GsgN9G8P9juC8Ob8t8HLrTs7xmgXedd9coolg8fo/ORF7v5fPDk4XbzjbT+0+JUP//Li9/+BP7TYu7a/2CVhyGKhnZ3zmAzbeeW9kGz3dXZ+jTflHRwcxFg5vH+QR9USKcDb84jwSp3X1ccA+/Efe+vi/s1nIIrxwK0+O69gvN9ffOyjv7D47//GX1n83n/q9y329m8sHnnkscX+jYcSTUP50Vt37j2xu7v3OKbLa4gye4K9y14H8SdwVjyOa+7h7Y3NPR4Lhce1Pez9XSzEw92dracxzn5x7ejsZ/7ad/zXP/NLP//epxIotuCRSiLSkL0ix3QYlN3xO9IzwEuzh7JONveJOVC5RoC5Ub+PWw27rgyvYSlN56gfXbpMfApjnwauKUZ9DCa4Jr8M59x3exuT1mM8M777Gq7Xiu2my/Wmm04+erw6K3GGI2Oo40F4LuAc/E1V3mOaRsNbt89655fbJKuRmcdoA+8YjhjfTlE5borf1ZRN8YlTGq5Jp9WISN54GqfZrbv3ojudr2xIFIdVsCi8Y6CtEytjcbIE7zCe06/TycNnCbtdMiRhhRmVlDPeBtuVvQ32ARuKkvZ01GFHpI8Y8mjicrGdELGztbixt0e/6xvDO+unHHrB27D0ho+Ri6vrFFNWN72Wei7sszxNwug4iAz0TXOgU7ctzjpO1Mtpik84D53E6i8XrEEv02Q7qfm5yMlFGRqv+Ewdodn1NPKxxBU6aLrpjXHCdVvnjWM61rYL/OhNGmMb3jxlnwO07+KItE0/apzzt9KbNPv8VPfhiTb1K8lmu51j4hCuabcMRrbpSDN3jbqWXR4tUx6jpk3HP+8Y1vGfdSl/PopZtMd5Spv6dbltEcXIPw6fqhcfrZmSWxzNh2VT0xWvkVuNP3X6cy0bepOXaYKz5XidkvKex20bTvKer5wT4vMx7OKrsOj8zo8tQ/5yiNmny4KX0LiJP3ra4pHLy+tIfOq2+XdUl809Vm3lCJS27eBiCuocAc8mDvrr1D1mX0m09sr6mCf9lTXfs7SzBmYNzBqYNTBrYNYAGvBm+AtLK0NJA1h0YtQo6pv04H8JmWGtFXGtFEwCbur5SyWW0fri2d/62OL7/+ePDqi1A6wKyheNkepsPmJRrKyy6gT7CEdIHQOCHFMszNbb6x1/vPjQB969+OD738X4seWKER0Yg0RGEG62uINMn1zf2Nohomz7zV/1NXt/7tu/Y/dNb/7K3Vu3bu2cHJ1u44S7ga3xeqIDHt9cP7//6sde9Q+3Nk4/9m/+iX/r2eeeeeoWFiA0fRlYXCnLgKGah5WSMCGBWaVVz6rN0qV2I+UOMWzQEwgSvhEI/BvQGypybjTYNKSWCYM0ETviHAZS5k9FMSBs0959GlQm633YFpxRbhnNbTi2AdYUcasEdmrcSa9xdjkNfDSN8DRoNs7mKTAaeuBJ1FvmvJxFPU7+HFeUVnjZfQcqrL9hCOvImfLQ45ufaT3lMRMVcWR0V+9lB1bWkAazcEarXE7y0ykrE+YyF+oDIx+/7+KAN0Dy4GL2y9Paj+zCGa0D3+I2ufuUFBJ9YsFmHWKhW+dXw3uumcJXimOeB2w6hRH3wD8GSDgOubyNMs5depiXs7WKwgs/DL22u7PYxphXA7bJzhp7D3ZkTiK3HDd4EYdw/Yiaesj8FvqSTZjUSwL7e9xYqNRLLvlOP/CVCr/l6JBcx4V/UzjXe9oERB+eqHHQ8MKQoj3gpU0qngevU12lFxTDaWHVso7EIKIe+RgzhRFOnJ4v6lj5uj/wzLN1/Z3Wm/c4lRBeHk1LvqJ4JBpXHCOkKnKq+HcGHOSZIV7Q13jXE/jFU6nOH9d5ovR8s8kkhWfG+zKSdvI43j0kK7XzpujzAuLgLrZ4RJ2C1wR1bn7qS3lJOWdhgefliSKr84n3G4c3fqQILdn2W0RZfKTSCE7ePpz9KnH7wEPpSvmiO/TKDxuh0/qTln3uQZak3PASWRKddjwcf0Mf9CXFoQXcaHbF5xrkWHCI/wwnXmRzwGijN2Wp9VUgvHDtUmavn72vGj8g8Y9eR/SfOHLpkDbySdrz30KiNJUDmMynvGc1oQOXHgTFTw2e+H0q8vIOaNBs4EhkmGM3cMjv8ZbpPcKz/RUJ+OglUg7JaZvTVdXA7CC7qjM7yzVrYNbArIFZA7MGZg18iTRQv4hLbGpw/CMQ964bWzhOLLch5mY8d++8dj4GEjZGrHDMDR0XZbAwJjfqlVMsowYr0HKFoK5eAAAgAElEQVRu30d/DIX8Mi4vGg3yV3lo0pobf1DUm+w1BjA2ggRQt5LBxNg4pnh8erJ+RwvyNz/6i4u/8Of/08Uf/df/ONFt+4uHrt/Ipv7gfXRj7fQJ5Dm49dmHn3rLX/lLZ8898wlonKKgs+z6D2PxkskPST5fYm+Ugf6S5gwYH3ZOAc6IbMOTsn7IQ6P8/M+2MTyTFIMvSivjUfXY1jpofVyuN6HMJVSE62SbRxmupc8e3zAxzBgSQw9HjuP70LFjOTAMCA3yMtpWczTF2X3ib/hypGjoleFuH0hjBKY8PoYOiCLZXNK0S5zNQ8PLV+O3bOq6eZdt737LEtXY9PG1xtH9PrkGVwF70EfjxToFyj2ZxIWhyjo7wtlw586dxdr2o+HfMyLRK7I2QSn8Cc6C7EPVRHSOwXPSkMVyyUA73SV/wTW69It/jImedMbRVjqrR1WNLOuUCDbeXInnJE2nPFZ549ruYn9HnfvIpboGB/y0fgSUlmS6reqFo8qDN3U/iNnuMeXPLh1qrXPrgbEwSY1zmot3Cts4pm3TMpcgBuQ/mC/0Icy0LoA6E+d0rQmzfCRTWSapx/umUnVXUzE9z/pcqbXWuM17rOi63LltkQ1yyRFi2mf/0oljhSTvK0lrvejg0wnUXDcOHTrK6LF0FsFT3hLpCNZjwfa1ABzIbrRUeEfQ7CfGlT5RYdRDfyAjShcnmpvx1wtIXH6h14zwNeHjobLsuahfzkuf5freWOnEcSVbtVmXB49yPBdu+Ys85nwvSMo2x/oYZdYCbY7zocTADsdZ8KkL+BE+sschO/hwYkmlg2BOHS6WNPVaGTmW6FF0vsULBiyfnxsRJ05eMgN+aenYD186sKmHHqNt87rg+efMeS3qPuGmiXZOa79yiVvb3NgjcHuPhvZwCuqA1vh06Fy+YhqYHWRXbEJncWYNzBqYNTBrYNbArIF/FA2sDNzPD/254Kr9i3y3DDpNn1XSNqFGexlT3PKPzuRpHw1YBe30Sgs385gDEwa73PkYdynThEgyE5Sj8Zp7HC+e+tgHF9/5HR/QOimoMjZeABonWmSA78G6zF94H5/1iNm2ZNNMjqRh4EEfbdIMiGGwrJ9trG8eYXUfYfoRsHAYhwFOA9yNxLQpxTCaZHNqQE1pCOcRQ4sOaWwOw6/3KhO+DavgteFzJA1Gk3A+QiWziYpJa300PfM+xN80hLK9U/OuHPUIUxmmRoyAXTGTJkOGvMWLBrv45MdID/8+V5rSLUNzZXgux2ABr3iqxSoTRtqoQPu0c5cTvRxYcmm0ujG3Tl4NfA1dHZw+UXz/3sHimMeE13ZcxzjPiCDTEaacNIicYUSa2GKUic35oG8Y6g23JOu4jB0t5VymbZxX8mIaWZWtaLiXEyVOOjvG/EZ+nINGs/iYnO7lJx57OI9ZLnhBq5E+0owO4Guq14o2iigh1X0VCVgOCju6PeVq8BMxm1FojFSw5fRoQXT+2L7EAx/yPZXTPs/+wI0850KcOGO8XhHHoYvGZa7Dy9zzZLlflegHW9KKngaPcp1xQcfYbtdR6nUMXHWtq7kf3bQ723aP+QIvLwyhZTh9KAav7cHhNLn2gQdl94nDVOJ4FigQ9Zwf6g748Lxa3zXC84d+/4ZMOm2cYzaFrPkQD8OX5wwDy6E9dABf6jm6HzzFfxplqb8xN8B4frgfn8l9xoyq0oGmHOLcGNcnI79gh3OIORhRZOXwY78v+POlF70GxJVN9KHNOxutDieUDuhac+J3nXM6JuWlGbRt8lYB1W0917TmH151wpscKy31vu4elfDmSzucpYRwKbtFMxojr3JCTM0k2cmFw3NKZ9yJ8vLTyil7n21usgZwCLppv49gNl3pGbEX3WS60bf80Z65EvFY98wUbVwzEMbrju4/Hrfn+4L1RwPn8M5TT31ih/M3bKupCHDxO7Z4nT+vnAZmB9mVm9JZoFkDswZmDcwamDUwa+D/hxrQ8ivr74HMD8OhDYjADOvlQlsPbviu/07yB46VGMYCz/lonhxrJmGhYctRx3qhwosBqOUZO4wU7zGFFZlRYyNEjdIXL5Xxsr52trG1fQRNg4zONHLaiRFjCeNK49GyhlIMt0QW1HDbTZ1bFkZY2zTckG+Zun2a29n1BpzisG/aH8eDBqRG4aB/GWYKP8VveydpGG8ljjy+5kRQTjRV8hXsZXzhIQ4nsDWYuBnXPDWdwlky2KZ+w6+qGcslfE3G6mzg9aIFN3R5GW/w6zSCrE6K7lfdB/eZTuTTqJXXY8tjHnQ0Sk/5O/VY+aezmp27TrY73j7H6QxrONrzBksfz6WtdEP4ZKLHgBs4m150GdQ4KIHZ2PYx0OMax/53N9g7cAOLfgtHARvigXLwOvTT8956bRY7t71pdVtoysdI1mF2pTP6qq0hFOXiurMnNBk3xbccN/Bbb/ql16Ir33VuSftiCs8uhqhVvnSQXIRrmoWzxqc84Kq9nFD2LvkapOB6Ka9Njaf5lb+UL+nJasNWvtKV9Wazyiuee0zPlzR1rLCALEYX6mOyDNM+5Ts8DX1Hp6w7KVhu/NlikpPAKDEVKD6dn+ztyPtMiJRiHR2SHx1VBFnzmccOYb4ccrzhESeVjiMdZ3luEFzZB0wAUtNzgOVjHD4nPhYK3USokcu7fTqePH0qL73arsOLSN3A6IBq+JzDY6xOTvbLrDXENYYIX8rI5rmuhK3wwZN19WG0m0eniq4ufeTrceBPJB/lGkcP9NTzdM2WrAWT6QKvMCZnQFh1U+8hgC++0hjD6Xy6gSNw901vetPem77ya7Y+8TG3OsgCytj54+prYHaQXf05niWcNTBrYNbArIFZA7MG/r+mgbbBJgbG75zFMtJW4y7XVz1fQKk5bRRaL9gR7IpDKiMkXRbbsnFM4Ebe9QBOP3rAtO3zlR8AX1YNm+oQUUGgARZODE9JYsRhnA3bMMaRBlUMVnJT19vhY5uCaEYFAoPOgu5Ac8zEMgyHoeb4TlHAqhqjtvEKZ7lplzG4AnasSfytxW5r/J2LK1EsDteSxuhzeN4eRzXRL1iExVrxK9Ipr+IKbyOCxPqUnlEXGuVFq3iLQSl/pCmu7MkUBdEuqEd4lGZFqLRQjU9cpuK1aNsitBFIoriPo8n95HQACu9jXrxmjh7gffIYGkuj2D3A3ENIK905oi+04nBwAP3Io1yOCyXndjg69NCd5S2ZZUA3f4EdcwPwMvlIcnQAqkSOEdlj3XE6xV71yA1ekMEJgVPD+hn5epxH8AaWU5xnRl3hyriod2hlHuRxyFBrqCJySl9iMBW98FENwV09Ogt0CBRf4hTO+dE5UNE5vUYYgfwNkxy4OFyZV3msGXG51bwNckvee6yPesqEcL410mSfKXzKE+2NTydlxgbC9V/yZxpHm1kwOA5+ooOB077INWhJsagVXfno/ubDMa4b6/TSD81iVc0s+XX91/qgP5zRB4Av9tDPcorDxyWpSqQT/DkBQiF0Q0MAB4Rn6OooIvlYZl0PXAOlBx9Tvs++e/cPTuIQu0cUpY5inVQbRFBWpKTzyvyM6LFcC6hvbrnvmI8aElmGPpQlOqckHx55CysdR4cn43FF3yiJg4+1P70++fbLbWgamaoeSheFTx3o+DYp9/IcTIsfzm+d9/bl8WsGrSfaq68HFbXmZUMe1+WNvDSDfE6i+qItfJMX3lrz8rw4oY/WU87FHRxwgjPIDxr9WE/kmXQd7fjMdWihMGB9myZ0ScyL6M7lhKjU09O9r/3af27/bT/2zu23/NXvWHzX3/jrgRfLnK6+Blwdc5o1MGtg1sCsgVkDswZmDcwa+FJqwHv/3LBPDYAvhIGLhusXgunSWC0ODwlodnQ0GA6pRGwZtXWEhWHkWDMhvLC2mVt/OVJZTWDe3Ng+OV9jr7Q1trKOURaj00csQ1cjq41YeE2bue0enbo8hWkjW5jub/iGazxdt386zrq8XIbr+pTPHmsuvj663jx0++V8Ctf4O5/2We5kv3jk2dS8ajQ3Pdu73DRt6zTtm5a739z2Hmtuvdvst82kL+neXV5MSi5PGswxc43wIsWRKJz4MOLb0TLFN8UL4owzDw3GdWqaIFvSN9JF2MyLY8d4cZp4eUVyHz92vEZ4nG+04ppaPPbQNd7GCa86+zLmoqNmOt+t8+ZdxE2n19A0D+EB07x3Ll7L4WmUp/gab/KlM6foLR/lG+MbT+NuutP6tGz/tN5lc4+m3Xg6b7hec8L1mIaZjp2WWy8NZ974pjgap/2WHedxOTlmqsPL/V13bOMx95gm8dhmrnOp+xvWB4Nrj63JXLPCZeng8HRx++7B4s7tg8W9+8eLI5xX9w4OFzrLfDNx4/Ixwy2ixba3cGbhIPJtlTrNpOdlb+rUclXqhPu/2Xu3HsuS7L7v5D2zqquq7z1NzgyHJCiZEmEKAvxmEIL1OQyQEGRakk3DgF/0YH8Ug/CDHmQLkCnIsA0ZMk1yJHIASpSHksz7SOTcp6uruirvedK/33/FOmdXTY+HHJDmdFZEzjl7R8SKdYvYZ3r9a0VsAThffBHg7fwS/heri3Nk+DZMkS+K9rs1Ut0d1/4QpPNzuH/gm5VXJ7yl1auy8+HMPbPG/AiwCYz1GWi+dfIYgK8e1fJLeLGlts8dVHbu8UOdoTaeWdoLQOzfJ31b9/2iAn+nek57bnoOaguu3CmAh366r2z0ZybbQnFtTSSAGS+kub5/fnl9/FN/7a+jwPjdKC7z+457YGaQ3fEJnuZND0wPTA9MD0wPTA98/3kg/2FuAGUwMLa7eG8h3PpjIErfHtz9eVrZccVChxcjxkXHn8LtknecRiaCQJxpbewWqmyIIWdDa7ynnh0UDZ03bd3uuO5LhoNR3WhzjgzAzOZwkrzPuJEJw8DQvvzV/FpG69F1z+GxJCb1isy0DH0N4CwNDHlfsoVj2FpFUCvPLchgQLcNzJXjx/GeDwaQKAsE1cVMGO+liA3QJoinLt/WH8UIpPVh+TE6JFvEullO2WEbWctxbWdJQ45ZO/DRIov3+2bshLe6rla8GTV9tnk4+a0+1w/U+V/siI1M0u4hfrBxU9SnaNKEfXZvssiwrpjQqFz9wAC3rPU9aV7YAx48gKboGxChZsMhXWorJiwZfwBg8dbrD1eoREIKQAOH9uvezVqJnALW5KlvBEbyhlWRQYq87RMISJ1L03p1npcFeCCDdmRE0RMv04Sf65Q/R5td2f4XkRA8UccUurSy3hEicTfXetB3pV/pr8LWLdrjuXJXZPkIeHR71iaMKgPrxXWVMfKET730oJ6rwil96hRQOjSttV7v3qeda2UJNlBYetr/gr4+t47hU9tApXOWyq/y9Xekfbh5iUne+soPDb4LP5TKFI3nH0goeuCCXOPF6I1P9I/PDX/DFOQVnVMhH8Gxs1O2Ul6s2U7JE0hmogCPc3FLluQeB9Sr1z4glQDYEWCUOjpvXs0cW9qDWmHsuWVuz1Tvy8vLbKeMPiFQi+U6ZOulGVp5twr6CbrBx/+fkly5e5xF5viTHY7p4tn0efZZcfnYrj6e6xXO6Gpb2mmoLMjSudptrLmMHciRn0WbpEneGc+Gv8fhnbk5iC+c9/yeQG8WbeZMf/LcHeRMO/SBp+OkzTl5Gb99cYljsCMn9JOnVzI5qJ9RRx9+4Iucy65eH87rLHfXAxMgu7tzOy2bHpgemB6YHpgemB74PvWA//2fbR0jcCB8GIFTBQbfp2p/N7X+3JQn8DGzzQj31gDOYCgBmREbzu635hmJ2Z5gmmsHYNYt9iXASs05qvYOrgSXmr99zYebDS9pl2VDs2wc963LEu7oNkla/ss8Wh9ppG+Z3ndpPn1tWnktQQrr/YFZhocPpr8s1/b0ba5oHhdVINt8sgUKTj2+dVBP790GZglYQF2fihDoe7cGmnz17NlpZlTQIXMSsMrwFVJdvNEb2UEy4QZfAZLO5lJGCrQWz1pyXD7IbR4M3I6JC4Yf0ad0QiD0AW9EMnhrZcvQnj3k3gBoIIDtXge82fUe/QAHI5CWpj/lE0W7FqNWvpZz2H6DKn2OtdjeZUtTLemDzOuSzt6ue21ezcersv0EQFVXXcRf67wFBoqXv1fNJ9eFXtW+1aFl2t56KFO/2taf7lvS2dbj+2r/dypNY3/zrevWB/bFVuRbSl7p0+Pt9777Xa/dV/TV1357mc6h0jtOer3Z46o+nnjorEviiwfOTi9XT588W51fCnk6rp7tPdBW/XV8fBgA9uBwj6sZWYK7ZpINYM5nx9871nN0AvT0HLPTUzLFLq5y3piPSp6nrK2yaw8gyXH9NkjHCnz5XBRt2AWg0i4Pt/eZ5Y7ssXqxwnpdZz/6/JodxlOeQb4QgDMrWVMCwXlw0y74uwOt9gMX5ypIXv6p9eh95gFXqLclda7yMkOt5kBZcBm//dKpd4F3299m2z3wXxCx5me7Bq0jD4xbenRar07uH98/FlAcxQmZ5RXwwATIXoFJniZOD0wPTA9MD0wPTA98f3kgwY9R0aIQKixq8/ZP4gECrTUBji+uTAYZlwRA7VFjK93dga68DYj8WKTv4n2PH0FTd+Vq3y5ZFQZmBoiWHuO9gZlZHi+PXfKUblnsy5lPquFnBIMbGgLJygx5UVffXqc8g88RchfIIYthmzxatpljEYG86A+NfUFEItT7EZQiM+eajfHyMaNowTZboRiQbCTbDX97HctXWbLVT9ajq/LgbWdtMwvVRl9pjO/dBtZFXd2fpU3xq76HLs+Rvoq/kKEks0bIHtkUxwYwgEjZFL2VW+wJb5W3AZ7VASfvaTc7rPSnK+ADctSDfkGyzDdb37q43cxtZju3lU1XmTVk1AjOiQNiOzk4uEB9Wx/Fbu8Jzik1o+E/1pOt7QPvHWNdqGKwsnlTyhy8BGvpes43BJlPbCGzyCwhMxmj04Je+U5XSrKsap6TTkRj5nn4QZroxADYhZdyu4R22NltS3twb9kHsKSu0nfp+77a3ry9hreiGIuTq6494TH6Bz/ptQsOfMqHXpWZdnUePCHIXNG94Zs29RNMIavMM+WkD7LL1fkTQKqtgY5Tjjpw68dqCr7P2kRPlodr/jnbK898eyvr/eiItXS8nzeiHh0drB4AvG5+wzJ3PlN7I1NPgEjG9fuDemyfvM6ZZucAZK43bfNlFJlB/GRdPT3Y3yJAmufBe9ouWXfrq8vVIZlr0h4dHGab5wH1+BUkQZDOQ/stWdHw9RxB7y0H+hEAD2+RWehzp80bB0Tefta7vqk5yIMC38ypbYzzrZmtt8+fJRmWrDUzNwUYyTOFd/1W1ry7HMrv8fP4vTTbNC/XoK9/R7TbLDL94bZV7D1CxMnx0YmS+PgU7CK6+NEwyx31wATI7ujETrOmB6YHpgemB6YHpgc+eR7oQO+Tovmfs75GSYmUCGaIXm54xSaBPgFOB9cViBFoGS0afS9KB19Fs+3YBFYEZfKxvz/LzCtH9FhCtDBwbLct+9M5vppG3hVEE9AZTo6xGY9Mi2DKkt+WxkBz2+c9hEW7MDPtQ274SUcx2LWvebSMuo4AOpQvftnfY+zZ8iifN/XLdO1H6VMMzgmU3dbWst2StQ9/d3c5VaenZJCNs77MNPGcL2NUQlsOK0I21YzNAWV4sAPqzDWdLWv4snXzGj3s183SCxo0ndfhm0yr9z2YPv+su6bMlLnmfKh9ALHrC85Mw577x6+tTgA2VreAEtl2VtG/ujoyY4du7af2S67QeW2/6Lsu7ceu93iEpcl57VLjBVBqHXf7y9eSrSO2pfXpddLZrq1Ty3PEto3WoXdfm2PTLPW3reV0u1rY1h9plnQt72X+zafldb3HNn/77SvQRB+X/l4DyvCdMVYpPb5q22/5lQzAIMHLAFPb56rnQZri4TLrMeiAvPKt9kVSDuX/6OlzrlcBmI54IYWZYq6l1x4cr+5x3lfzLWDZ57T4uP2xl4nXS7ZqnnvG2PPLtNf7J5AFUCUPz5uLH7hXv/ZPr03bfLulD2K2ZvLCjAMyxW545eMewNkOWyvX68qsklZMMu2AVDdkV9JS/tHXPpc8o8qAIf+r34qSW/prR/rzm8D8D2N627S/DbDiUxlt5bOaS/lpix9Br/Irft8d4PVoi++gucK/PrfWdb0yzDyNHfzeyDu67ewcs0X6tcdPPrwH4en20a1nTZ1nuZsemADZ3ZzXadX0wPTA9MD0wPTA9MAn0AP+R/4nqXy/6Lu+vfZwfiMwYisvuU3wmsCI6MaDpzuTw0wPgyCLV+3w2vcBYshKyJY9+uTm+80a0IIwY82KSJTFRTkJ0kZwF4Lx1bw3gejg1XUjzI1sxhT3Ghx77DcK9bAiSuurXtJWqGxPmdj98qxSAWRlYdAy2rvft0I6RnMsvmkvfiNgLb3KXzmjy35wmBpbGrQ8N7kWcIUvkEHYXnzDlT5l9D2qMSsVoOqzAXDFF1SfPwNwSqAtCMGWRoJXeRsQs5GWmwps5SjQJuvoJLoGkGbJWW7yjtwQpN3tWAWYYh/gWAXkKqQ9lAEc+IZA77uEtQjesCPzD9iQrVxuK7u4XL337ttkY7FmOPOp7HX88J/szBhSFDzMduGup3X41D6BwwrTkiUDzcbHctMPlGCDzmVMw5Zqriv8/bPUHNYaV5eaoxpXOm7BqprXwQj/h7m61l13fNu19CuwImNC4TOh/NJfwFONdrs+uJg96Xg/te7qKnhR+m1tcEjbU8+2/hq2sTD73ucGN6K3oApWW2+6ITe+QKE14+QpZOKUhz9rqPzcz4C6RDo0+qvk5rkf680MvNSRG4fBMzbk3SbS1wzlHEDGu5R38cn6Zo/1/jzbil1L+2yfPLl3uLrP5yEvfPA+WYKwzW8GfJSjnn7yG4H2V2yjPAMYe/6MLZWgYrEZe7x6PlnOLPPxGXqmv4yC38j8gk4nSMPPKr879ft341tleW7MNvN59IB+ddC3R8dHSK85MENN0HDNP1fUvDoJ+CuZcnp845r0l+5i1M5drUOBPOW7Vdurz7PnDVpSp0ngTVDO8fb508jPGPUC3dGMfzIZ62L8Djm/ObcQOfrN+cpcOxYe4Jxqirj49PDq+ubRaw8fPUR50Hp/NNQ+5bs9Dk03r59AD0yA7BM4aVPl6YHpgemB6YHpgemB6YHpgXigIk5DqBww5S4eA7gEUrc5C8dAjwAogRVDvBJb5VrBEZ2jNM2ynjbCpgSiBoGj0/qydKBnW/c59mUZyzEJpqGpIK+CXoPLDn57vGFbaMbg5mm/oJ2lZX7cPWSbkrGjFts2PVseZgyVjPZbMegXSrReHfA3C8folWRlcC8Q0KVlSXNNUGsxaG9ePSZbEek206PLHmARr01NsK4v/BDDGvZyi64E94JZZpikSEMJb9bD5uwx1dEZdhvZj5ID8hNMD3tDgy2OXToP+mor/mJl+v8GXTvr5eGD+2zRIhPlHH0MqQcwo6jeJuu9fGVd9pecllXrwnUAoKS6S3u411dVtnb2mhkdY4wyag3WfFonswYeoR+reSNjw7f1Km5LHkt7Wi+pvLfPItjycol8GuXln6XsLB2tN7/2g22Wri/1WLa37B6fZ0UR6OQY68pq/ZpOHt4336bretP1ONstfU2Fr+ZhXdqXx22zV7d+if/ViTm4Aoz/4IMP2Vp5meymQ7LGPNvrAWvp/gngWNY388j6TkYWbDIeUEdd1qBD52QyPufNr2dspzzlzZSCw9JY9jkXz62/pVeth7ahbfNqW/2ebM+k80UBgmQe8O9PzTWgmc/Z7e0Ztnow/3G2eLrm9zm8f58tztGNdRagbPgsWXtuSdVHwH3ZhonvladX1O16/AOAfF1D+1n/2/UBy/hX/rF7rLe2pX597CtbbK//D6g6UqJbz5H98vJ3Dfk7t/4gqR98+RcXt1i+A807dD5myfY+6qhLXz+EDpnlDnlgAmR3aDKnKdMD0wPTA9MD0wPTA9MDn2QPJDrBgD9p5GFAZXzlqc/LbW2VkVDBsQGYAVFdK4jtegeS1v1UxFaBcPe1XwVmIErVBCAD0S4BtxgcmtGovA5Cm87sKrMXRjwWnaQD+UjA2HqkjUHWExR6uFFKeco2D8X2vCB7CiqrYFOy5tP3G4CLhuJdgaYha8uSlvA7fOEQuQae8sqZZIhe+iQH5G9mrPSS1jtPx6pgtHSRs3L0mDQ3A0wwMy0HhdN+AHppnHwBWABxfOKY/qBF4Q1mnETvykqqzBCDedrdU2ZhnHLURBUNxZU5Uq9UIponU0ydke181nzRlxQigbLS13lN0tfgbUbKjeedIVPwwq12b7/9JugemS8AnUTc2Mr8Q5+10WBm9Hat6f9Sr/1f+ioAmWYxeoMd6tR+d8tpSgMnGzslxebqZWytTe2zXV3KC7gVJwfHEnRhRM4fizJl68bftjG2dZC3fKInzV6zNrm2DZIv26mlrmZq0HRtq3XvvdZ64TrqTTtM2tBZ73GOEWjpDKToN2TK10/NaenFQG+gKB7yiRyVs+AY5ZuhZ+k14XPQRZ71/L387Git60+bBv24MqTkuEYFZfCkIOjzZ09Xj598FD3V44Dn+f69Y0At3gCJLm4x9NxDU9qUyf8ouznM38P3L849iP989dHT09Xl9VVs9Ry8k5MDACIyowShUCW+RZfaoome8BPkNfVKe/z9CUCd9akPlKPONbZ+ZzmYH54X/Oaa7XbDVkzH3CeL7N7JMVsx0T+6mrXmP1YUiJdnbLhDfp3JJX/feakQXzaQ7Dyeo8wXD07Wgf5CPw/l9yxCwbVMXnTDnuFXaWKHTCk+j1c8n/tcq710cRpLB8dWn/L29333LCLIBgUuO8Rv737wwQfvIOwP8PcCIPOJnuWuemACZHd1Zqdd0wPTA9MD0wPTA9MD0wN32wPEkm7eqmCFAIgko9sbA0gDQgOeDnW0NaYAACAASURBVJb6fhPId+Q7/CNdfwxQLV57fF+774XAmCiyQm0CK4P0AWI1rWNb7hAXvkv+TYvGCfakyzgCTK/dvxzf9/K2REd0XvJdju32puvxfbW97eq21nu4pJtHEC2OUGf2dAcsSo9u4Bq5Hc1ST+A72u1LcAsIUCAUW7NM/6NkS9eI0EMDc3WM/n1lqkKft/Chzwikw8Av1oBoQnTgPuCY7RqksstCm/4PKuDakcZAn5I5te4nDTE0tpjdkxVIuhi3vMHyfnQMGNd6MmapW8AC2mQXe3KfSiCYBofabdJow7LYJjDhmmu6pom9wz7vu30jK1LgFoAOW0qRAr4WYppeua1DPUtbTeTdcwqj0AnaWmxv2da9l0/z7b6X27rdMcvycnvr1O3N1zG2NTCIBzZsah5KL2nyGc9Q89mMx47iM9aez/rwqzRtX+vRfbAddGVv840sO4fcXhNPnz6rZ4qF7ll7h6xngeKtqFrD0jvf8rkChD07vWJb5vnqyYdPAcZuAMrIHKPv4Gh/dXh8wJoru3t+HB/bmjHzb18Belt7QhSQr+6EUN26WGttnezO2xtsO7hdnTUvfvciTlCYFwr4Rsxt0W/+lm3XkWA+yWjR162ReU4F71zOglbY4bZLde5sM5/NrY+3c2pbz4EymyZbn/UVPymxHUGZC9p6LqT1BEv6d3yebHdrKdNwfHt4+6n/+Kd+6v2/8BN/5d5vffFffATnUk4hs9xZDyxX7p01cho2PTA9MD0wPTA9MD0wPfC9eKD/I/p7GftnOeb7Va/v1WZDHfMp/qSlA6Hhj2uCHDAQ8xEM+QxuK8C13wBp6bce29dln9k0bgO0rftbN9ssfU3gNToTbNLtmB7ntQPUQZbMsc4es6/7m5dj9EfzSGBoNtGQbaDmLSEnABOBKYybX42RtkCKlhlbBNz45H6hl3U/6tH3jquzvQqwqvrWrtT18rDVoDaeJwhtvWhCXvlDekv4qzEd2qjNLce+fYABElNyyDiIlkmBqzUNL+smraXeylcyWpcc6L+wv0DLKCIKkHH5gvemPsAElCFIH7l43FfBP/5tqvBSPrxu0E25ZqncB5h47803mS70ZW48Q8mruksj3nabbMfyt215ByW8vJdni7Cu70QdtDX9VNNuHx8Bi1476tY0DsuHce0n7fA+vNAn2z1FJvj0uNBEAedEDrWOWqbb7Aq8QBbdyiyfuKYKuGkZXgsjKX9bD/9xTWXx1WtfupqiAd4MW9tOdVnKkIW66Oe+onWyEPVd2hljcVxspT3mjWvzbpq+Nr1jeg6973n1CSxdHbHgLxhEdpa0kVfdlYm2mWH13slZe48fPwnolCwstleumZNTzhK7vuAtlKeXq/OzywBi+jOYLbzPTq9XX/vqB/l8+OQ5B/KfR0cP9jf7bN/nimMZb0isFWAyk0oASH0ueDPl2cX56vzqbHXN21b1UWzCKU0r4ObH3wvb9Ffb45MbH5M9dgkod3l+zmH+l3nDpVswe53oPwFkPIPv60wys8pqXbD1E3u8z3wyRct/t/CcOn/Dun8jG54q4wsDzIJMMtnws3PU8+QWbbPbaptzbQ11C+el7fjhZo3dPqd8bEfvnauri50LXrYx+BxxfffHf/wnPvVP/ukv3vuZn/0vaqGNk+nGlM7LHfQAS3KW6YHpgemB6YHpgemB6YHpgY/zQAc3+Q94/8P8+6Soj6Wv3ydq/bHVeFlvwqeM7esfm5GRlzAL3wSE4Fq3Hta/Gd5BlQ0dOC3ntAlts7+L9+rY4z+OZ/NZjlva1fde+775e+3xy3416HqP6etybN/Lo/ubX/d5ta9put9rf9qurvdY683X69JG+5als0+6/eNkLun7vumWvO2Tj9kxBKtWCIR9W16BgC3DbWc582ucwSSvtsVr6NSTdnnk6vxad33YRnHcx625jJc26E+tC9v6UwAaPjog2Dfgl10yaG5Xr90/KX8BkrRObauBeesnr8hfoAKR23opf1GktTQv71/2Xfc1H2mW98u6Y7tPgMRPy5DuZV5Nu+ThvaXHSbOk6772w1bf7TMaBnwtxza/Hmd9ed98mm7Jw/vmJV1nBXW7V8HzrKHFOrB9Wdo/4cXcWpa2tYxub3r1XOrXevs7JZjjy0JabzPtnjx5svra176WNfTmWw9XDx/d49yxI7Yp+uyS0SSISxFIBWJaXV3erj58/Hz1lS9/Y/XNr324ego45psmd8g685yxyjBzQIFFAldmUvkRNDo9PwuY5b1t5SPO0EOWz7J1NDWDig/gGGDaxv/wlL+H4wva13O5Dp+bq2uAsguAbYA3wL2rgKm1pkqnmkP9Ufxq3fjikAL3C4zdxUn9DxvaHV8iSzDd0nPQfGxdzoXz7ZiMoy9gGG1LH3hvu9cG9s7Oz3e437Xt7OxMsO+Q+jtPn370/sXV7aO/9p/8dSdhllfAA3OL5SswydPE6YHpgemB6YHpgemB790D/sd3BzTfO5c/3ZG9RWvEd3+6zP9/4NZBzp9UVMcnFTJuw5U60J2oiKjNc3J6zqQ3EBIT8dwdPxVMbSU7t61PB1UGbP3GR/ttX66Bpu+rh8SbdWbY3/xeHqPE5uG48K3GGJI26sO2AiysQ2v2RuhHoO7WKe0yS8Ri+B6d0TWBa7ZnVQBrk+uk9BIfckwDgLWlSAbpD+0S5KCBYvYHXxlX9fJZ22+mjoDVLtur8oY+6JXuOi1b26riN9KOwtPsrryRjgBf2n0DcPdZpZBKxnxmTlf2o4cfSyZ18MOANfoBSVVgrMOcjaVYm0qp8pEVeERvwQhnYQBuskdY1Izfsa/b4gernpcE+JDxjPUsqcO9dUAKs8TW+GAHQEF/V5aZ6/AgbGy3BADRVmXZEB9bLcXLd0N26M2oEXirdV1ZXo5zRukb47bzK1NLjQsciIw+g6r6FBvHZOkw+60G1xfBHtn7lHXpbES3ueonZ92/KOR36NEM/9nfdgt2OJcuq9g6+sUKy/YSEt8vBGpv7OcweOk8PytrU+up+8x65X+bUuu9+UqfnL3oJuDkWss8qC99VZQvk7HWrLFOtTf6kcFlYdVFH+8z1t8X/pqP+vZ96LElWX+OBfQxM9LD+R8//tbq05/+9Opzn/4BwCe3T5KVRV/rDtaEfA7iP2MbJYfw/7t//9XV17/xmC2V16s9zil78OgB52eZ1UUmFHNxyRsnffasW645X16963eSc/7IMqs53+M3hO2QpKWpl/LU1/Xr/dH+UfmGta5r9MY+c6WOzpW/Qc5xxrKMPffM8f72CTR5vpd61W9TzzdMbmql8GvNc1LzJU3OOBMIhOe1k5h1qQUlqzxO+8jOs51aSv/e1vxv/8Ej9mRNmHFZ83Z5UceJ+fZe+30JiNfLy9Rvte/2YP/gyfXl6/dODt87OTl65/T09JAFAFqvdouHYMifl7vjgQmQ3Z25nJZMD0wPTA9MD0wPTA/8GXkgQdGfEe/vle0yCPxeeXy/jEtQadC8CXf+ZJp53g0B3Q1BzjrZCgafBGkGoRUgGfgUz6oblHVo9aIs+y19la4D1SWl/VLarywFNM/lWO9tT2AsHaX7UxlfTdeympfg01B9Q27fks5+6xlD33KE7dFvM/rbb8ST4ntc0nKXMhxhfbhmQ2N75Ornj3Hn1s7q7CDWcZbwJDhX3/QBknlFZcAPwDGKW0jdJxW9ogPKMiYcrRO8W6yHBl246QZAmOGXUMHPOn8bf41x5ufcONbi+Bg76ou28mfpZnNAGcbdACrcf3iyuufB6mxbc75vAFUCIsBLX/gRBOhS/nFNbNeOfbGDq8CFqliktV3/+PG+6UrdWiVFV+rbr746w/nR7pK5lTGYj0vxaL42Si+YUi8sUCdtKLoAFtyXDGrOlV0qZOE++nArz6XsyAjYWbT6yYylZVmOsb3AMOQM+83GskiXdbPxY62n7vPasutautRLKyqrTxpL9ELveuuiduPv2LNdR9L0+lGuIFDpUDxcEy3Pdu/99Llc3svSN0R+4xvf5PON1V/4sR9N9tg1mZM7ADbytJiJdcVWS7cufsRB/t/65oerb37jw9X5eOPlyb3D1RFny7uZch++zgnTHP19q2TLltfxUW3JBfAJmHXAYfTaoSxB9wPWbPRkjl2/BV7Th5vTjn9dC/s+s9qEHK/6QFDJte04TrfPXDZAfgOSKZ166Y96NkY25QBXbbeYxeZa04cCfFlT/kBRlBPQL88pPh//YJDfL+ibh7Te90fZgqDX+Dv/XyEwBy9/R7xe3l5g/z7v6EDvvb3ba7eWgm6eHOw+uLpev/9wb++zJycn78L2K/Dy30JKIcxXlPJmuTsemADZ3ZnLacn0wPTA9MD0wPTA9MAr4gH+A/1OFc0hnPmuNn08heCXAetKgIwEigJTODdnxwCw62YzEHslIEzWDwMSJBm4USrgHWCFhKNUcFWShXJSCCb7asYU4ZwRWZqW9DYYpNmmHuHOfYX1RFdjjCOVb8CZoG/BXx7Ns6/NMwfJw2+X4E8wxiymZHNRL9oKKgNwwLvf2Ka305+MmEjwa+hqYK6mVfQRqo0ygJzhM9/c2GctxX5tDaBXAI5kle1YAIJ15Vq0QZvlf0tShgf+W6w/e/7R6ikHj5sp4tlWmQ7s2/Elc1EPY5QzFEsm1QiWw0SHWpAVXzFHcTUZI+libALvBNrogkxn3EynEOpHBvinvvGfI3GL9gie5CD6DtAB88j7Wb3z5qdWD04AHa54pSrBuNIy3hWiHQIFsBnxfq0/DDKzSrf4Kb8MPzOPgkDqbDvf0LCWXG+gFuJU1mlVXdYBflbJ0abeFtet4/ciXDWUWXNif+kDM/nyUZ+SV3LjB10fYCEjIrf04cFDZvQI4GV/6UVrdIfjdq5VFP167tTON37mTLQaSn+tvyW4qT7DHKgqo0k+0RO58QvzCGPsu2pOXPXBsNVnjJq0cQVndEXv+BErM76GOMq5jp8y79XON2XMv56HV525xX2AI2dDEgeVrFuFKXN8pNg/OFx94+tfX33pS19im+VjDtU/BLQCpt055JwstvjxNkqzJS85R+v584vVs4/O2Vr50eqjj55nvh49ur+6/9oJb6o8XL324N7q+P5xnlMP+Pfcr7ZL/8R3Q7bPXBYya9/fi+qvbYlHyqf/8LCexX1+P+sMMQ1yNskgw787gGG+RAAvZLyAl0UQyvPKzMxTvvzzfNOeK89EnnlfOEy/606fOdrfL9erdOOx5B6eqevvkpVnlfUSefbZTkV+KJCrgGZspt2rRblmp+7wDAr4+fzrCecmLwMwS87nJ/LIb+Q3iWf2iOHvXl5c/8i9e/c+Dflj+D13mCz5WEpA3c/vO+CBWv13wJBpwvTA9MD0wPTA9MD0wPTA9MAr6AHCk2ztIcYiprlKoIQbCIh22OaTWFWvJFAyiBr3HTh1PR3jyz75JIjj3gDQQKxLj13SdQC3pGld7Ov7l/tbRnjRGTqDR+S+LMexTd/8vBrgfZx+S9rO5rBtCY7Isy0zu6L4bIPK4lEUtjZPdTPjp/Wmg3t4GbAKCIwi/TaTr2zKmLS35Io1DbndIrYmkPZML0NPt+8l/G5/KMSPgXpkcm/ozv02VBU0JNh2utVHEor0KYNFxtgQGhrdy4YvaRgsxzxkUH0ZQDfgsbt3gH7nqrK65dy0R4AUBRWUrMyfoJt8F6XtFzSLvwzW8b3tARCQ0aVAg63uy3mWxjFy3/gC1EEszrJpG2ZXKybqeyq9BVBgo+S2nn3tEeVD/Rg3N4KRbuA6EIeyaQBRgVIKFJavxX7LZg5SK+CiupQxaPBZ7KJefKveZmR5DRrZ9Li+16/aVGNLtyEuF8cL5FpKn+0asa1l2idwU2qVDj1mSdNt4RvcpOavbW0fWPejlaUz/AdodM1Ze7bdDDDJN1JeXHBmGAf0nz7noH7qguzHAGmeVfbo0WurN958BJi1y5ZJM8GG3jA3C8siPRbmvnWxIpAKlIUuPCOsvTUyD1j32VrJmlbDbI1kHe0GvPXlGTxTrG4zCMsOaMbcinQJzLqteNf7mN9z55o2m1J5W128FxT1ap+/sd57te4jcIB+gTpZb3nGdJwsxhj19+M61nfJ+nOyArDSN57G8EVDwTEz3RxzxJs2sW51hA2qu7tPHTl7ewfgtWTjuTUUY/m8TvcPwv89rr/FR4DMUsbU/fy+Qx6YANkdmsxpyvTA9MD0wPTA9MD0wPTAq+ABAx4DorpiMXEgZ+kY5ySDrEEEA1ODHQM07w3irgUjGO9YQmiGCPRUhgJM0242k5lhVPhfg0ZbzxJfRT6MclWXLst79VBOZEOjnC62d1ne27axTZBoBPJpGwOkL5ot+BCwajFWmQaZyeBCvQSPHp9jMIlowsmtnGF3+6356zvvt5rCR58OuwxES4/KFDEtR9rakqb7tnq2TbYZnLvtSu0D0kS/QnU8aHyfk35KFybWLYkE8EbdsUkJCtEv+t/LCJAzZ84FAEDAMchQQiFc0XXMaXXKZOgoQ/RBQGR5CH+2FGZ+iy60gAPaIW3ersnB5AJ5ZkDdcpj5mw8fAjTAxpOK4BlaBup77fGcNPVxrF5Vd/3Bd2gr4wb+XYZ9VuMPM+pMfyEDx7r+SJEHPM3EE2BwnXeRP5IDZiqni9mLmJOMH5trfqo3LuTLdS6AsgE8h7z2t9w22iqHuVKnAkgA4tRFPq419RvUvS5a//LBoFVoc81YqtgtOJM1XCqWvT74KcO/ApGMV2ayCodf4wP8daBu9DX/5JM5F8ONm62j0UERzAt/pS/DsLHG1/3Wjq1fs0aR5RrssbKLjc5ThqIvwNg+vzOHh8ex78MPnuSAe/V3bn32nnz4bPXs2Sl8yORi6+6nAMQevf4AcOw+2yoFeOr5O7+84Hwxzl5kLTp2n5dHWNRV0NnVuPa3hKIel9DohjVbCy3+LHg+2cHYKiqfHbddQuu2zSw51vy+Z4x5JUstmaKMiz8Uh69cmYJtvCklemi/JRoIOA3/Z41kHtKNnJp7hGbcIbYJqsv7ED/Endxb9+3CaB//tL011/FG6aNM9B7TWFlvJaq2rmowZX+fY8XgeYPuWYvYrd9PTo53zJ47Oj6Q/h7ufOPx48cPHZKB9aVZxWjROG8/+R5YTvIn35ppwfTA9MD0wPTA9MD0wPTA9MCd90CCMqxcXgmI3GLJ5rbaBnS1vgED4FhtgjI/BkwddBmyBXCQmCIf+/ueyqaeRr7SP8KhDW13cm1d7CtQbkTdi74mb3BDWse1fEETSwK71gmZDaTYu6SXtkC3Ukw75S0oFvuEaWJX9de9QX8i2m+zUX7LIn3GMLzv5et926tMwY9lmzy6/+V7x/tnKX0Hb+qOsd/zlny7XLLItIeg1WKGi8E+wnKV3nODdkTD4iR5mtUlsCcYIrA25DRqI6OPLWWrQX3prh8LtIsPGGP2mKXr2QJI3aQz37b55huP4tkOzKXTngYUuy7w4P3mbKbBU7nFu9bBFmisteQsxn/wLDoaRmneaQcA8OqneQoqwD76LccoyY+8LWV73Tvec7qQlvbuk8+y2G5T1oL3VKIHbRmDgMz1GGhb6WaWlzqVn4s/fdGy5rzottLimWFXt+oTS60n7wf/ao6BrZt08mz9in/5s+7LOHkKvDTQ1h7qcfJpO5rnBnCDf5eW67geqwTBw11AGAGy4+PXcuC+b281c8kFJVD87FkBZO9+6r3Ve++9s3rzzdcDjO3yMggBrX4Lo+urZrF8ECyMZ1LZl9AFrMPR/i75jwI3bEHVvthLiyBawEzYqPpe1g+H92dWnY1MoIs8z1sAWKbH9V88HFfPrnYLAOub7fotezcynXTpECadeqYg98AXWQAuWvSi/Tf8HjjWNew/cDjadoFTeWhX5NHjfElr8Tm0XzwsVxr8mRBKi//ZAprxY8zegS8VABJ0DEvSzGTm4+DwcO/owYMHhxCLes5yxz0wAbI7PsHTvOmB6YHpgemB6YHpgemBO+eBBDkGUAZYq9Xp6TOCrJUH9F/5L/9X54ArFIOhzVkz0BkoOapLB07dZMBnMdjy04FbgjHb+Rg80VsZFASCFvvDlYyfDgJtD60KjtI8bV8W62nbkqbbtgI2hj6t6BhstKa8HJyuTiMw3ATlAxRSXwsWoasZdFs7pVWb2IhDKrhFd4akHZ6ht56MIILP9JXv5aw5jq/QtcfSbwDLHyHu8EXZ2YCa0IiBNQKiobcG69dkqVzkTXPKgq8A2a3gmLooZ1u0P+eXwcMOZTlGvVJQLrZRqfmNR8tO5UKon5PhRGXHt2nKSKNG2fCybmXblbFm5+wAxr3/3lvJysqB5edLLV2H8PajLPnAI3PufQAhfYNks9OG7GTpcF/nMzHA9eUB4vhVfh6sbrkGMNFvB+huSSv9rbfPgb5t2d3uNtS0cc04afiTfjmf8Z+gBb7e+FI7JOwij6H3ZusdfXmGEL4EAzfrc2QOabd8sxYYk+d2gB/FVoiu4Jr4KrQq6XpW99Lf+3wyrwt+Ua3WnuqKc8RSBEW2HJg/Rtg8dKl5Kv84Kl0lD70dZ58ZU0BdQ2619da+rDRkJfNNnf29QDfdJADjb9WOIA1vi1wDxj4/u1g9uH8U8Ebeh2Qw7V3srt5688Hq/U+xttgeqK2np2era84mk79ZbvrkBvCqM6o8E801I3Ak3c26tmcKCsk3/vJZH37J8qOVFzemX3Cu/EojJXZA63PhT4z2eAaZ7ZZb1qy8USa/i05J/fQUReraH9mOH/f40WK7a4INnOjEPXZuzjZkQnARKtZv1gF8WBopez6rYd7/MACAxtszC9g02+yKUYNYOY7lKoiuTHvU2yw5X4yQttIlGWTOj7+tR0f7t5/59GehdrSfWe6yByZAdpdnd9o2PTA9MD0wPTA9MD0wPXCHPbAJ4si4IB5ccyj/FQGPSErSAIQItsF4BWGdXeDYDtg2fBjYQVL36b4lj273Kv+uh8cAzBzTcnqsbdJmHLJflpk6geWSvgPQlmE8WuMJQNV/AHryTn3Egs1bWoPkCqyjwUbf5hk9oeti8CnYYkvxXPQZHS9K93vN/QAmmqRlFLdqlU4boxv+MuzNeOeKeSTzL9kx6p2CzAETJsCV1iIPmOTTbeIetznvSz0Jvgdt+iHNWVtaNuYpYKA6a1dYjXvBA7fZRhJfypEXV+6QQSYN98mQYewuOrsW3n7rddYhb8QDNNE+5epfA3Dv2x+ytb5s857W0DRdy+/6ck15/8J47HC9BPQY/JXTY71/udjXMiI/Jpau0qZfPQNWjbrtC0ZFU9lIi+YXdGtdu791KpvLF85nz7n0TeM1Xke3pY+87/HNt+t15l231jXrhdvma6v3ASQBQdxe6fjuZ0opWZ0vyJGPoHu8INATb5S+TmGPd7QlOmkDH8daz7ZnlyeOPDg+Wj149DpvqyRBi7Vr9mSeQYCbt95+k/PG3uCssQcAr6wliM7YTsmh8eEjkNwvCDCjTIDMq+DY1WVtTdSnyaSMNtecVwYMxT5gwSIBMX8bPNjfx+noyLdbAg8EAAR4xZ7AxQJf6G+pOdrjbDCy3QbQHnCMPnllrfAcS69PfTKcTz+b4nMaZ9VvQXzqnEMgKBUZAT/rd1TRvSbiP9Z6+7L0qgy4NSD64e7hRtZu1i064Q+LPHzDZuviM2yJLlzlxf0t2zh5lK73eYfD6vDg8JyuUxx2xnX8KHE3y531wATI7uzUTsOmB6YHpgemB6YHpgemB+6oBwjcUiq+Wf3e7/3B6sd+/K8S1qxv+Bf/G94Gt395c52XAxoEmVllLHRrxGOgSeDbmQWyqGwcglfBEupmllmWgZvBk+ADEVQFiwZ4qW4DdeOqBFkwrcCtgq++9yqNZdnWAZrZJQHFhl0h5Mt+6b3WfQXahImxx77wHrSeLWUxAN/l7WxYmHpda2z6m+841PqaQNJzgizqEd8NubZZ3+pQMm1PEgt9ZZrGl54CAWVnAwPlM7dEqhFDGFvKtn36/PT0NJ8KR5FpgAvzyB6mxI8E5AJZjfJU1kozfimWjXLoVeLgVfprenZ00a5s38KXhkEXvTTSAiDg6hFNECRL3/DJPk5/cP/EKUy7QJ86qrOGtn1hM8Z0m1c/ENpNGVcBRAN6YQb5ULxWRpnz1Oui5LCpmCwyM63K78UTdeGH5RsefRZe/Dl45tD6IUM5KSI10W34Pj4zW4cz0OiSb+Zho+5YM7TnWUEPZWzfllj6OkZft/3KCh+u8QUAI+riS+AZfMAo1UhJlhmmhwcaCBK5Wj1HyrnVS1BHbt5ciyLKkmZvx7OtnD/1oI3JNztSf7IZW+fSr2Dmd6xhWMUHL/hKn8iSImt1SzafTqHc5nmSvf6QlzTVV3aHLG+tPD4+5myvI57Tg9Xz0wvOv+Ienp4jdgRYJWiliY+f1Bss85ZICORnttQaUM3tyAWMCZgBzmZBa3H5wXmqTCgAMACyoyPO+WMrZ3yNLzpTKucYouYlb9D00P49/YEf9uMS7OCaLaDamMek57P8oFVmxiVbknHK9F8ufBPmZYA6Z0c3y4t7AK1kwFEXZPOZ1A6B/6wx/Od8SetV93ofvZ0Dc84YV/Nb2WCZX2RIs68yykMPeauPPmv6ANzwk6d8lE1hKnbpAjzc27tBlcdHBztf3rm9/iaLq1KTpdK9s9xJD0yA7E5O6zRqemB6YHpgemB6YHpgeuAV8QBB0K/8X7+4+smf/I/We0fH1wY1HUAZtCagwhVe+argysCRYKu2E3bQZqC0DWT1nmM6uK7x1R+eI+BNu6gIRdgtAR336tDjm15eCfQI9uy3ZDxX2w3SLEs675s2nXw1P4Ph3QR/30nvGvGiHtop4FD62Zc/roJjaTewV1e287VOclJH+1uf1qOkbPWy3dIy+rqkU9ZN03GfQlBu0GrAH1Bs+CixKDoRcyMEHaQ3oO4t4l5A6wAAIABJREFUeswnRjX7F6+hx8KKrsvfZsgsqKIfXtC+ZUfbSceCum61UVDsGjBkJ4jqevXgwQkx/1n4BGgh8M8WPmjjq8Gl/dZ+aubtJ/XQ/70ObO8+39DoIf329VlzAweIDM9oAjccdpaVsYtRgjXy0cfD46krv0CJF0FFn5Gljn0vkEyHw1LkaanvGhMwNXDVi+tGHqX7do04bsOb/uYXpuOrx2UNIik0sIg9yhdTY2x/bPceysGhQBllB2Rr5kN3qz1WUE46LbLN0jpFd6GnMc4MNIEX9doT0FvQ95syw4Cv8I+x5Sv96HT6HF957h4f31x5yFspzSSzCOgI3FxeXq/OzslOjP6ll+2eWxZQCX3ye0A/6uSeCQ/4dXx4tDq5dxSwzTfe9pp03fh8C0YJWrkNVj8qQ7nZsgtYecKh+bd72BlUUL+8OEflN/jCQ60dHz1xHa20cdg+7fyjRXzQIFXPUeY0/iy/3iC7eJb90ksj6Nylshorc4w3T8YmrwHlhg7yUIYArTrrH8HAzqjrfmngD1afdbWGZs8tpLjvOVlyXwKn/M2vfvWrv8dKNousi6b24uq2eb0DHpgA2R2YxGnC9MD0wPTA9MD0wPTA9MCr5YER3hsgEwT9j//Df7/6/Oc/f/vzf+/v3+ztn9yw1ZKAB/yLjDGBijXn8BgMeQC0wa/ogHWDeEtnRgU2kSeAh/2Ej0VnICutIM0YU/3QUpcyddlJO+pN21eDPEvGKH/EVwIRBpRdmnf6kWm/xUuNLT4G2IJMDffIQaDDcQaDOwTDFnnLM3rpmAEs2a5OGa8dCIp/IIyuBInuWNRk5QpQhY8NYVy2b+xBnGchFYizpW17vEYX/HtN9ogZIMrh8Dj0JkhF5z0yWzx/7MYsIg/lJyj2fC+6Vze8KZIIN3YoXhI79I+2mriT88qcEdv0nTrDN0Y4aJRsc4MoujsvCiDAT8mFLxir743nn8V+7R1rgHp8PHz41uuvsx2LIQAWL87zYAm9wNRmHlSMovxNUT7tnBM+6ATDWL+AXo7L/Aj4KRvjnY+Mz7wBhuBHVS/bvJaufdVMxfmpFRTiiA8giQ/qwPfiq4qtc4iEOpTJx2fGPuVbdyud80kvbaUzdzWsv5kPdXS+uqibWUoh9QI/LvFhsq+GjF7DNS5Wok35QrBEm9tO8Upt7OzEWiDlD8enD77213qhjTE+kQWqd8Ye/dBv9IVeADKgEuN5qqAnnMaxrV/84Zqk3+LV58s/+cR0nit71cNxfgSBTk8vV/eOOf9L3RmHdRzef5G+a9aV6812wTOvDTi5zpUrQNfZgccnh6v793nbJdli9454UyYPh5ib4+SjDfrM+31ROvqcT9cu6sDvdnV+dZ4st7NLMsqwybdcWsjQDd0eQB6Dor9XH0dnT56Cbz5PyuEJir3+/mqnnlOWY6I3pKGgbUd0j2K74GN9fHEH49DxCt7q6O/Sxud42O2dZhwqV5kCYeHNvanEnU2mr+o3zXVa2Wfaq18ogmSwit7+Y8uX+f+Cf4Uav/78o49+n35N1DKL9xmUWr7KP3HmtnHefcI8MAGyT9iETXWnB6YHpgemB6YHpgemB6YH4gFDJGI8wY/b1R/9wW+vv/6Nr16994M/emWwQ3Cz0wElQY+BDDstK6B2288yw8VAyo/jlleDWsdU7FSggJJHMBVaZQSc+Zjx0rZMg7Ye14Fdh1fKlM5in/e93ck2QZmMcStYK2MHRb7LOC36DzuX9khrn8WDxRvESgNf0sq6aLzXF9Xe19a3x3htffpadg45w6amj27w1T7tkV+3RR4nHlk3g8yAOApoC3S+eY8Q3QhWqcWS+2STWZOvY6J3zWV0or4p3vuRh/Ipm17aooPzBFpQYw3EoRBoRI+wYqg6rgEMPDMtIB2R+/37r7EljiwZQD3XRGaTAeEDR+WEvzpzLw/puli3hLc2L+q1DbDAEfWJ/9w6G4W2fOVvUx1CX+upZTZvrw3ANEDbMtWx5UrXAFjxtffb9bPPIjCjxNBuvTrsqeeq1718W6+lvG6TX7f3mGWf/V3v56bom68+4pkZQHBoAWv6pQe61jaL45rHaEqbM6avi67mpultS/tolof1vgoy9/3y6viMiyB4MN4ti66DZIzRcMoLRrJ+WEf9HIytf9FTkJTlkecjgCS8BHC16er6NKDYG49eWz169Gi1J2Ib5Kuy0ASYtEmdlCGYpD5jZ2jaS19BKP0HTwFfXgKx5nkJrWuZdrdgCtoJaEchjaOonzIdX3Bt+djfBc8Eu91DHorIK76A+oq6YCNPVOwQpFSP7W9m1dUFxSNDcK/PYuMFxivfX0zy8Gbc7u51xkeuv6mH9TviVlrBOPm7tspeNddE8nFpZz2sufw+3b+En37x+bPz3/r5n/95mWNgaOfXHfbABMju8ORO06YHpgemB6YHpgemB6YH7qYHKvg3FBthLuHNNfjI9SVB16VBEW9uI7lsJ+ev51ymEZAZAPWnA2OvBksvF0JPgmpbK5jqgE6Iw/sel2yIMXhDgxzvlWXxvvu6PbFkdZZOGGMmT2e2NZ1ARkF8xVN9YAcowR03e4AlobURwDB8tRPeARi0zzEErgFPlAOyU8GsPFTQD371amScop/jhWTBNL3nM8WH0Cql7Tdwt73tXNo+GJae0MR35Vy6tj5C+OrZR88LIFOPpAMhSH0joOZefsn001/YHx2cQ/0s8OQ4iz7xQ4kU/YL+BumCa8WTHmnINFlQUi+9ULbuw1+aQSUv2sy6ev3RAzR3GZaemQ9lSsO15kd5jEY32zI3Q7f0k/EY+uEX5yj+bL9GHdci800aTKvXfl6bQpexZkvWVrLqq7XdZ2OpftY7ulg810rwaHdk0AELpn355XxFF/StLWv2AkhS0DJrtnBoGmDrmtrYjU7aJxBT9gDO6EsIY4M+ob/5OzD94wEpG/AtHQFEWePmSd4wzjO41N/xfizKyd3Q2WXk6nfthxf0AchH/0YuEmTh1l1lWbqvdWg9ox9rL4YiINv2BOHGpIQuK8L1Vs9En8WWrYysgavri9XZxXmehQLJBFf3V8/I3PLNk+urAskEhy2Hh8cBtq44pP/58zOyywr4Msvq5N7B6rOf/fTq3bff4K2XD0N/zoH+As01d2Ymkk3ls4Ev1A/zAyL171hvPfTMMD2mx+2DKmv8Ep35mQ3IdksWmdsmtf+WuTTDzBcGbOwXDBu/E54zJpjnnCSLl/eoqIWcrwN4cc/VuTTzC/QtejnHB9k+WX6teWEQrwi4vZY/aw/95KGetdXS56OeG/9/IJlkgHmX0B9xzpsvF3Abpnpe+bKNm11+ArK9kncXeO7b3u3B4cGX+IX6Rbz1jz569vSf/9zf+dkP/89/8r8pmALzDaRYLfP7bnlgAmR3az6nNdMD0wPTA9MD0wPTA9MDr54Hksaza5x4RbBzBRBgNgARuIFSBcYGUH4MjAJAjYDaegd1S8cZQMrCq8WxFmmbz8eNCxFfPa7H9NV2xzV/25u2+9wGZBAraLHsk3ZZuk99vDfrLPoJeCDDUmd5ca3qZnjokBMbF7bJp/n2NXxo98B4+bX+hr1dbFPkckyPaxqvoVuMaxrBtwYGBQtgVB90W5s9tnNEbKqAkqFkZQl6JNuFuVoLWDjOEptYAioFDYqnuYDB2taW7XXppyv6l7/LPugjT0nVnyv8txlC6qOuN6vX7p0QeCte+QKS0AFY7RD0D9wpw8PbvqGnV4P42AzFsn27/sY6GPMso6jNl/Slb/nCPsfVenVNlP5Fs1gXjpN4UeQV+WJXFMeol21bXepZsN5yi7ra3Z5me/N23VlfFsd2Uc8622qr99Kmli198/Gag/XHVDcv26X38zJ96y9N87Gtn50ekzYGW3dt1XXr5x5begsOF6jWOlBjcNXQJDittC2r5Qvs2K5/z84uVseH97heJSPr6uqCNYFugFtg/mlzPd3nHDHXyh5vnXzywRMyqMiiItvyEeDsW+++xRo8Wh0eSel2TDKocLMvbujfQJezMyOgVC8VGHairrq4btWvXgLhOLcnUm8AEjyUAx5XB9CWv3ZX+9wfkjrJDy/zWPS6v/0U/43fsZ4DXhHgL/PqiswvgW3lxW/wCKAXBwKp+dxS5CXY5QsZtF9dC6wXZCyQVvBRX5b+BcAqW357HCKm7Gve7LmLPw4OeFkDGsiLcsuVf2dQD7Pldv4A2n96sLfzj06ff/Qr/9nf+JkPfun/+F9ZnCqtZSixmWGHz3LXPDABsrs2o9Oe6YHpgemB6YHpgemB6YFXxAMjDm1reVnZzvXh/j4x0c3t5fqSQKreNJgA1UBRBIPS4wyaUifuSSBHILYstnV/aM10ITjr4E8AJeMI9rw2j753bNN2n/W+r6C0gIHIQR0l9jYo3qUGZ9qMbL0OfVRTPn2ovnAMXDd8m9ZWZfhGvBrb1+K3w7k9ZrPIftOfwaVTB5wQEVBKUwEoN6G/NZMpOmmT4TXt0GW73fCTelZASx9MEvOW+A1ol7PSNEp/cnn65EP3dsHJ+aHBrCzOQVodEpsypwb+xOLwq6wUprYkD/+UQYY5ar0tlS3mYHSy2fmP4vg5c4ksmWuF+lhk3nTdRrN2m6m2T9+abWM/8rkfUjXItZMP15yBNmj1wWbudZIFfq4r+7K+NhlIpXd4QOMbMwUE2o+qoZ+iexjVl28HDRiSWVCemXXOR+nb22qlybzJGz1dJw7pzCu0SrvYH6cxASUUCKGU0mnb75bXBnIFxzY6wxKzAub4HFpaftPEtYxJxhr0AjGqIogTn3CmlD6rsVzR0bHXKmZ1+NE2i2NSmEt5W+JzaJWhLaORDgGqsKSp5jx+zTg8wHVIzrljrYfjW38ReecNOMpWZG4YDr2FqvBvFr3Psvo5556jB0i7QwYTOj15/GR1fXYLwHUfkOyEbLBDdNtZ3T85WL319sPVG6+/xhtS7+WQfeUHJIuv2dILQLbH2V6XZKNd88y49dBSWVKesaUvzbTz7ZQXAZqOBLpdA5DqM+1oH6I4fcNy+orfWJ/wFRAkTTcyLrwCju3waAo6uX3S9a9P9L9rFCm5r7XvmqxtpZDAbPt7FHBKN1rQK7890AiMiTDL8whA6xKfOW9uq1yztfTw8BAQTKCwsuy0w18r50LgzbJDJt4++vl76UsKgNXkd3txfUVCIvlmPMe+kICXI3yZ6i8j8xceP/7WL//sz/z0B1/4wq+oM2lm13n5yzA9fOfX3fTABMju5rxOq6YHpgemB6YHpgemB6YHXgUPVKRWlpoJ4PljZpGlnYA9mQFuxdsJolCBn+QVsNXwZfDbTlu2Le+736vB2CawHB0GnNL3GK/SdH1537wcQ2C20alpe+xyTNGWHbb7yRZSmNWZWCU/vDFPHmZphCdX5YwYOiBAguHRr9taZuskH99wl6g19/qs6Ja2qkeXj7uP/KhtYC6oIpehn/YnDhY82M1b+VYeyH/A4eKCcvwJOqEI2TQVvhjUrnY4Y0n/KngEw9alyycKESQLqFRUvbFPurZVsug8lkeANPSwhMax1mOj2SxksbidjOB9fQFvXirw1hsPIsbwO3+o4NgABeiv/+IDecqYsqmr86iX78Z80WZdnyivildBD4DClwGk0Nd6S4aQlPAW5Kgr/lPnAVgVvxe/pXt5XnuslMt79TKrZzfPlp2CcXpgABxsj7t2bh04ivbIw4/+TD3gZNnX7U2f+mbsAsgJVwGc9kuPKJ+5ZjI2SFmtq/oNGP09CQxb8nCMLJdyq63moaUEHEsF+6AvHiVnyU+SHu9VyObWbY8seDPUBJZEMZ8+fcrnGfX91f3Xjt1luHrjzddX77z9+ur1h7wd1TU8/LW+4U2p8uW5FM8VtNoF8DsACHepOn8+s867QJmA2hUg0dEuLwAYD3/WsCuV5+Z2bNH2+e/+gGqiailknakzvtQGn7iAY/TtXRfoGNsAvHxMDnk+ekkMBvBdzC+Nrh2B22Rz3Ra4dTPWpfrf3ODLWOnvWr0ddBcAbt+5OTqq89nUL5ljAbwCqkUOOtTvQ8lRB8HDa3Xnc8TZbPiFn758drNdef/2D6n+8vHR4T9++uE3P/8zP/2ffvDFL/wzhK0P8L3u1juymuWOe2ACZHd8gqd50wPTA9MD0wPTA9MD0wN30QMGNwRzizA3hyxfHewfXu3sXIAJbUAGzvGvQHx3HOK83PO2DNxk5qcAoS3rgDnys58Aq0sytAxaaVq229/y+2pbwBKBHiJDA8RkScAvGWNDXwEGciPCzzOWzM5x66FBY3hw31u/rAt4dGZXcEHVc5x03BrSea8evYUxoZ5GISffm2i2/GS7hSF8DFQdr5EVILrV0i1igjDqXiGyZtEPWW1/8lr0sdvhCLsi1ow+Y+oMOsF5ihZ6z1syqCeqjx2lB4EwTeoV8EZdAACSuURrsmQkMK2MbDOYcY/9nukFXQ7vp+74mltuJSPglm5TPMNrBMGl4/BHssqkK/oAENrPWN/KeAHoYHaLbrPPTBVVMPC+Ifgvto53TvhjXOZT4Jb7yGKA+UaVjcVY6kBxuUarAWyoq32CY30v32WJa3F2AzdLsCxyIY5cFI75+LPkFZ+NTsMfgpNZq2Hoimn9K7On59lrZGO76xumG82sJ7uONoVK2+tRgMdiW7dnvHRK82sU27OX2gxDMxhdVKNfkdoXDTHFXCKzt7IsWQee3WZrbB6DtDXrh3FlF8xgkDmhSX1gGl1r6zNt9uMLxeaZc6SNDFxf045sn4t9/UUJmIqcPq8umuUZXa1e5+2n+vbykiwoDqFXrm+ffOPR0ereIed8keV5zZbLuJM1G+AnXMM5+u0AElkq+RGZmKnaAoLyU8cD+agbMxIfo67PdSHTpaeZaGZl6WNfDKCsa94AHBBU37EezD7M3CDPM8dOz89Xx8cA2WQZHnLGl3IvAPMO4muGRH6/NVPfq0/51cxReR0CCgrA+RbKm3rVZp6d9QCAGcE4VOX3xixE3hlAwWbqZtCtfVEA1rRv5KUc9aYxW1QdgTTbby/YhL93vbsDOCcVOPzhYzKPf50ssv/l4vT5L/2t//xvfOOL//IL/qDB9HZkjpWP5DPL3fZAPU1328Zp3fTA9MD0wPTA9MD0wPTA9MAd80AC1xdtWnN2D2jE7RVBF7kMdQizgRIFchMGBC62QXsPHzSppp+gLdcam/um7av9fpbF4FxeS372S2cgmDOyRr2BCvs39ASyQDg0jADSTkrz7THyI/8kgb9g1wahKvINP+nkvbwOkgTHxpn2RaDf0JasbrdNorLpZT7W8xlju96HkdNcPAfC0ePbXkV7H98gx8PBBfzOzs4CSiR4J8jdIeBOBs2wRQAKQnxl0GxwrA2LAp+kydHcPrNXWa6B9qf60LAdSH1nBPY56F8QSv6DRoDD7DKH7QIm7Dlf1wJgN6vXX7tPX23VuiH7LbwHZ+9Lz2pQvnUBMfu63n7x+vJ4Rwq62N503vspFWvNyncDRLlGovuL/olsxi2BYuGDpdzm3fI2Y4ZN1i2OEZhw3ixN7/1Wz2pfTpN0ebGCdAKiFNvCR90+rgDQIAo2tU6u8f+S1PGWtsP5Kn80s/bduKJ7rY+t/Ng51mvzWdrmQ1czh8cUN3gIxAlERQfa2l/tJzUQuHG7tM+4XLTk5OQoWWNnZ89JRDwL8ObWyocP7q3eJivx8Mi1sF0n8lGGn9bvdoBaAoeI5jmqudg16xCf1Rso9VnZKUDlllMBWLXpt026VVRgS777+0fIqHUYEAp5gmfqIjDWRRrtErAinzDzJ4h2DegpHzFo11avkdK9RrcNZrhZwofbPJ9o1nY6dulHl97x4Xb7rWN3Lj1vbB1gz/mSR/PvezNsKaURaJv/HwHfJ2Qa/+t7945/+YOvf/Wf/9x/+be+/Jv/8lclOyi0zsdua68MZrnbHpgA2d2e32nd9MD0wPTA9MD0wPTA9MAd9sBI0QhUsr69uDgne8z9OkQ0BqJGggRnBlQJsMjyMETcBpYdMJeLcgi9wdDInDHaNNjKIdLw2id47GBJHspIEMbwDsbk1MFgAj3oWp70FnUp3VINoKFs34CYIm+KNNI6vu+9GtZabPdjZkXkJ4ul2tNvlkvsCfmWj0BhfFbtrY/Br2f0eP6RcWTrbTifYjMfA/zu60PglXOTgBoadIxcbqPX0F/dZdGZQ1rbdPq59FitvvaVr5BqRtBNECz/nCVERou4RfwEH2X4p+1RShVthz7qchWwwqkbXQNt6A9KsrVumU/HGDjbjv9wQRLRwseFk2IfHzPUuAYoI2g3oD9Axglb2z79qXfYOue5SAIIXLk3o06woIZVdlD8gc6dqROfqPMo7a9Uk7HDnWaoJ8V+VeEuH/3mFltLDjUPL2QK1sDWebJ41X+Or1koP2Uec8uYUPpVsnrsUifBkY1boLRPHSxNnwpfATVHe3iMgd471zghpNrjWM+BChgCkBO+kmB3ssTk43wJ0oQ3PGKPUE+tc8f4gTL8Wx+BId3gAe1eBbJcGtLJO2OYE/nZD3XaemuyS0ya9I3xUISun4V6E2hg6+I31qLjfKYsVwi9JYsrvxswy6+R84QFuuPe/SMO3L+/eufd11fvvfVwdXKkPy7QF+iJc+iSwQa/gFuM1w5tLD4xKHJcc9EXnursM6RbfNtktrxyLXvMqZKm7FX7PIPhgpo8D/4UHBycZF64y/WKTLcCxQoE814eV/Gf+jAOgW699a2RFvnu0iad+lm0nGpKzVHxNzvVdaCl12Sc7rM1tNZ//Rb2eN44GX76Tv7yPgdbD8CObP0j+OYLC+z35QSuVaA1Hvv1zs4BKcg7t3/EGY2/+uU/+sNf+7m//Te/+rv/9v+OZlD4TypOfCno99AVxb5DqefmO3TO5k+IByZA9gmZqKnm9MD0wPTA9MD0wPTA9MD0wP+nB/yX/nMyNM7JEiK6EhjL2TXEhZXlYlDoJ0EgQZjXZTEIqwCuI6EKjKWR1rFdpDMI7LYEYASKXpe03S99F9use/UjfQWAFazSGVKBGEvr1bxsa362daBs+8eVpSzvm37Jo3nX1SD2Rf3ka9Bqu/p26XFdX45r/gblXZa+UY+ABdhgMXi17fnz59QYI9hEhhYRPnX0EQoZtGau7GRr1XaOAmwYkKseQXxQEOjl3npxWyXt9MhPYJJzmEC+JKSf+cHG0mrQp517rmbeCKJ6KL1zc48tYg/IIFvfnAbEUJZb8EDf0p+Mtw2bMbfQ6E9t9tN2tc96TXS99C/gsdsc46e28+kx9I7Stb6GyND0mGVbZxrV9OhfIceyuvSpNdBjdOxOwOOtz3stSK8vlnVllt5bnsu2eFr/Q2fpdT6qqW9ll8yMZwakZeCmu/QtGu9bj5YnYevi1eJaq9VRfVkLtDcvMxq7CMpkTszW8k8/+BsTPtwDguWlCOXMHra5qm/4wtOd4ZeANle8VVGg9MH9Q7Hg1V/6i59b/Yc/+R+s3nnnPmChaweQmHE9Nvq7vnFZ2S/70lHeG/uwy9YGkrZAJWeesdZcLztuX1yOYYDbRJ2pBr13ee6EPvW0Z5a5Xi3aqS98w2aXgMVHZnW6ZqQpHaPTAMSSszZk1jilVZEuB+jzzAvs2qN+rrmc98Y/TuiPkr0Yw9bRQ4C7Lvrl6orD/Nl66Vi3ivpYo/st88ljvbtzyW+KYCwyPwRk+zdnz599/r/+r/7OF3/33/4mPzw3CNRDpMNFfnOe11fFAxMge1Vmeto5PTA9MD0wPTA9MD0wPXC3PLCNrmLXLmfF7D7nHJvnBD7EQwWmVLCbw5iLSuCDwMcAr/oM5gr0sW6A1YGx7U3j4B7n2ASLI4C23fqSvsdJ22NzgDm0/klr8arMrocPgV3q0Hr107LDSxynQsjwSJu0o2ZAXPxqrECNfcmIkIbxCUAHX0Ng1ewtVdULHZFxxsE7w4Yt3rd93R4bRvuSd/Q24qUYaGccwa52Zg7oQo30ysP2c4PbEvwiUEU2yfqGt/YBZq0BJMxESwZQtpJlQNG77ZG/ZIcFhNtYpCBiYDWxAEAIbAADSLvj2z4DwkWh0iF01msOVFbfC46ywgI4HJLhIlZ3azAuGID/k+UH7RIcuyF7SJsbENsfAJ+8lmVIZyxnQqEXCqe75pTa2L5W2/oKlLoRrGFgNOXGt/gJgqCoiEfmuzrN8Kk16Fxk3kaGk2poHQNCwWTBY9hNq9lEeaOqAEx8v5eMpGEGfLHazB1Gu5VVX2T+4Zl5Vz/Gdem7onOxVYvr0LL0iuNd4c73ejxr12krGa2n/m0ZXrtdfmaNqdct4Fb46Rro1Vc/+HxKrzuib+woXYon80d/PUe2l13Nw5Z912b4MU/oCXFljqGrdaYlwNgFoOzVOeftoctf/ss/snr//U+t/upf+YlkkfmGRtejmU8oBn5bQFTWjnMDEG+mYkqc5BpWm5o9twfn2Uorj7ud+pQb7ar5KlskoSl6ab9z7Hz0+WDSByRzHQKu6QfP9jKbdn//OJlk5UvsQwavhIRMv9ePTHT2ee8D+FFFD2WeoJffeoCuGFvPBqL8qdlk1CYTtn4ja62oo+O0q+4FvNb767zVcn1c8ynu7bx6BiHyeGvluXrsmFXG2y/P2U76pR/53A//xs/+zZ/+zd/64r/6Vp6z9W29yWBnKIyITYmvN7V5c0c9MAGyOzqx06zpgemB6YHpgemB6YHpgVfAA8uQ5Rrg4RkB0TPCq2sDsAEsEL9VEK0/vK++Cqy6LUABQZd9dZaP0VfRV3BsLFbizJYInZElZdM/6rYVnwrE7fejbEvf97jlNbpB23S5WYwpPQ1k0RUyA/ZBPsJjg8KyVyCm+bTsriuzbe4+r362+m1BxKbp8X3tMdaXNMt7+yxtp3K73ge0p4Ev7a/sD1vwn1kjvn2Pw/vdLulB6/KWV/TsgUTLad9GKyHBAAAgAElEQVTo7zjXgLM2lolgEf2WZIihh6BOACqdab+udxglWyM9NByZy3E3RN4hI0NRXQ/v7bEdjoywi5oPk8fCEzSkdQ0/dLbefu9r+2VJGwX40h+CXbkKXGj36Gz6AsxctwNgaBvL1FA3rVcZyM914nVBtqH1RtrQp/Xbv3oei6bApdgk6Iie+v7lIm1ssL/1DG1Rti+sFW3Nt/eSt0yvY3jopF+O3ciwg2LmUbRBrHAxsxCgS9zIjviXdpdMebh8XmNLZ7MG7Q34uXuUZWJ2ZAPLeFNy+NW87yLzBjDJLcIBx1BYbPb09Hz17Ox0dXN5FRDox//Sj6w+99nPcB6Zz7Q7xAX3XZuMG2CrYGwXQaIu2hmfL3yoLZb29eYeXeocrvrtsN1tkHkW5KkfHMd4wVcbfGmENlvMl/NNkD4OwlxmwFlqu2XNzc2QrV7K8hqgEB5ucQwnM0LxW+YEn9SLKcom6QtARuoAbvEmtLW+nXNpej14rZcv1Bsx7bu6uMzbMW8AFpUtgEm7h1AqhCq2rW8+4OUCv/67v/X/fOF//4V/8IcrwDWI6fYHx3me5VX1wATIXtWZn3ZPD0wPTA9MD0wPTA9MD9wtD3B0zdrssWSQGTSOwLHOmyFwshhAWTqotN5t6eCr6x1g9rXHiUx1YN1jmp916ZdlMz7BZvUro9ub3lEVkA4awsmmkZ/3Ab2I73yzoPW1oMkAOgwkLQaAHSSnIQEmdg+9pFJfS/P3agise3pLFuE5I2n3lQd0JNODTKUEt9CaiWPx2/HFI0356sPiHRt7h84jwq45GAG422F9i90pWVjPnn44uBavjDWoNcAGYRDSuSKO5V10CbjVPDRcowO6NIbQtgh64M36EyzRfiYxftDoMTZgQSyShgwe5eoDAnR9urGRvjWH8QuqPWR7JTu9AD8AQDxjahR1svQVNKLqwduEaaofphvetmzoh39jmzYNfjJR71t8wZv4MgFrgLw6P85MKOyEVmt7jFfHlA01b0iKPv2lz2pdu8Cs1DVeoypAEvsZ5jVvLc1gfTTGYmPhEDUHAi11PheAiTPgGuAv5/0xJrZFHZhib/s3azjydXH5TV/bf8322WSyKZN6eHD1frvuy7asA3SQJj5Atv/brvUaL10fYi8u43qss7tYc26/dQT6yMM3l+YNs4wxC9AVKb1vodTWaw6M94UcOXMMm684T08Qye1+57xHxDOyPMReyO6dd99YfeYHP7U6OT5gm6VgLesKADbrM1LrS9naF3uRq74+79a7uB7ii2Gr/i5b8T3PmX1VxxaM9OkRfNUXkuZ3DX7hIT0UVbRPWQBs2NtnMh56ryzGuLZc0RZBKTPMZBt9ocl6df4yIbTzLLlCnS+zDmtd0qJ8P/Bxjq2rheMtAocyrnG2wNsW+OyzfkgQWx0eHwWIvMDX+9h55fltLkoWEl+Z5v29nS+/+85bX/j7f+8f/wbOfkbOMbxvFCu7MoSbWV49D0yA7NWb82nx9MD0wPTA9MD0wPTA9MBd8MA2MixrfHvlR9zyWXNYfwWEhEQ5g6wNNkRaFusJHEdj1SvgSlA36Jd0Buw9ptuXdVkZsFXmRDG23vy8d1wXxy7r0oWGgNK+5m27n7SNwdU3AucR1smrebSM1jN1RDtuKdP2bqstbhWQ2i7dZnsmQahblwxawR1StKTHVkuNYWDZ4Xg+0vgxSK/ckzE+/LknIBZEOD09pRIlZYwtUEOTcQSyytY/lvgVYOCFQj3yEuvSM+S3DuGlHsTBAQGInXcAPbaAg7IN9wmV2kZ4ZGsfXY7XDoESgY633ngkqxRxgRtPK6fE1sV1Iz+92/62RfqXaSS1rYv3DRiZYdPznHbWRmXflH6bcWP4hv+GZyktnX3Rd8G/jBc42NrjfdNnQgav4g2YNGxQX8EwbfPT42xvmuZj3WfFc9vaF9W3fU6s6+TwYZ1Yck+74y191QeMhFcgoPT5tZ3fanK82+0C1QD+OH4PpDNjmUdH+7bS1ktsR5qcg+VzCKWAmKhixgqcgana5Lz4QgPXruCYmYa8QyTgmICNKM1nPvMDq3feemN1xAFk+4JBZEnW1srSZQ2dGaKu7rJ/XIfNWm17/yYEEBugku2eG2afJfOA/pkLbPP8vOw5pa9sGmtvMV+OrD7l+EGCzwNXs7I8QN/SMvzdCLiFzsp3rKXvU7cJJsJp+te+bVnOo0959TV/6eThmOaZe+i86u/8A8Kgc25tF1yknU2TvKUTQJnn9uJgZ/Wlf/f7v/Nv/ud/+D99ZbXr78XNIcM0iBkcgrmZ5dXzwATIXr05nxZPD0wPTA9MD0wPTA9MD9wRDxCBb4uBzVM/BEXsfCqQxADJs5ism0RQ9QEGQJyAC7gmgXnSZ6ot9IO7zRlHQCd9EoEUTXsHbF67eJ+Af7RZ7yDvZXr5drEvAexos9700nQ9Ydzoy1iBkgSCA6BQlaFOjU/obBAYHo6JPTEBXaOCA/QDQFF810EuETFBt22CP5bo6A06lF+K3z5Bc8bSbsl5TehVYXTRGF9jVXwI9JJ7evAX5zEd3ePlldf1Fro2QPohx7SQ/cFb/rb31XOXUCb1/mrfDlcEsEkGi0oYnge4cRx2CNCQwVNLQENpK4RA9SgE2hzGb7aec4srAcLYwsVB5e+8/RZQiUABgIb24qvE2gAB8c9Cz8yh7Cj29Xz3fdZhdW/6rDouWUDM9Q6ZSmsUFbgR9CkF4YXOkY36rPSMd47Ek+Qv5dJnsZH2bdYiRsWSoq/D0bFsuDUZSlDIs0rZJ6BkixpsiNUMuvhTGdz3KMeqz+YqMAYw1RT6IOvIDMaakI3+jlF8+ode1cZoZfCJPuM+xOhiNuQOmZAwKhqRHhViPkkoBPBhPTiGfrOO/NRbQfWjMkvYRgYZYwJE6rwfIEotmA9AGHW7JqPPtz1eXFzkzC6B34uLUylWrz+6t/r0D3xq9SbAqrsN9Zrr/9J1Fb/4O6Vq5Vc5pwhQ8WfWKKsw69n2ZJHCxz5NkqN6qkf8oRDG7KCnVri6/S0Q5LK4riwBwBinjmYjuv0yc5Fu2tGneXof3gE141ZF0FY8XZdN4wIULN1BD+2SnS8qSOHitJQOavdiKRm1HtRH+TLwatZetl7mB0x+ZXePKX2Sn7Zzc73eBRhDBV7gcrP+8sPXH/7+3/1vfu5r/+LXfgUe6JOnJBlkLyowa6+cB2oFv3JmT4OnB6YHpgemB6YHpgemB6YHPuEeMJpaRlQcf7ObLZYEZtcN5hAsgX34gssK2LS5gzzvN0GclVEShHFvoNXjOjOn+7pdmi62WZp/1/vadD2m6bpduoAvg0/z6v6+Ot6P4x0jaFPZLtsAsce2vtZ7XN97XRZ5CfJE3yUw0foQoJs9Yn9oxuDlvU1LmfY16NN22+a9V2k7VrZutk3Gcy9gR6XAK4N4xC95tw+ihvPghyKQZWl5LSt1aSIfG7C1aXps+gAOBM/CI6tsLDMAEeW7PdAiIAiit3rnzTc4oL9CbG1Ay/Bd2qmcjayM3q4vq93nmOJRtva49qFX16LtTTfYveAbQdzub57NS/pu67F91T6Bt6aVbnnfPJu++7qeLKJhq30fJ+fbxwz/wqTHeE1x25w6uS12+KZ12NBAaJt1/VNXZ4EVRHuXZb/0Tp+ZXGYCeu92yWOyuWwLGEmbwNjL4Jh8ihdjyVKyVDYfeoDeuLXPdXx+fl7bKrmenT3HjuvVu2+/sfqLP/bDq7fefAhAhV0AVbdkijWwVlsIS2Nl9HmC2rW17cXnXJCoPuXvjc08M/KIfuMaFGusz25ve8pOvbb1Z9Fs13TWng9iwDP5C25t12TLq3FjDqks2+1zzHI+neNl3XtLtznee8c1rVd/L5tOGus5hP9ov7LF9vdx6XrNOLqjz3O89TsffOsbv/3PfvkXn+ztOb9yYHJqyViZ5RX2wMwge4Unf5o+PTA9MD0wPTA9MD0wPXAHPGB4kwiOOMjMsWyRMXjyY0BlYOS9gdAIklLXduvd1vUQUqkx9BNo9r00Zkck64aAzaDN8R3QNb+ud1DXvJf0aJZ4VeVbh+5fytls6ayYcUurQaM4bgtOFOGG5yAL79CPIHjYvs16Kj3ExuCGzcUc63JTMra8rVs62PXA8mW973tLIGH14LT1uxzWZIDsH5jRtZfssQS9zJslCSmAFLdXnIC/fwQDM4EIlDMQArNqtM955j5AQ1K/lrZAkDmKYdDWvMVKl4vZQvwJRgjEbIqMBeYwaznHggRE3AnG1e+dt98M2KFOvnmwM+fKO8Utvo+ita56XbYPm7/XnjevvYZ7/ZkV4/wIYmV3H3PQfcoLP/yZM54YH7na0H3eVLWwEqtDDtZj71Y/7Xa87bkqF9pKC3Ng+dEXRli021Igj5lco16X9KXfbK7QDg+1o2iL/gPAMffH7E/PvyIDKPbK1Ufc8bGNa/HasB99NXW2ui5S3DYLfa1XDnUHEBMUKryTrDH8ZLJVstawW/2LtvQ1a88lH49AlwwsFoDcr1k7Zok9efJRtlOeAZJdCpAB2Fxcna8OWd8/9JnPrD713jvcj98TxviSiryoAiZmSKFt+PoMZF4z2cLfnlhWjvIpyxsjAxryG+ccyYvh6ouHYi61WivoSHfsdI2PaRnrCJuyxRB7eQ4iR374orZLyoX78Tyq041Owo95yQNXs81c9wLGzokauE5922UBaj5XLhvnruZgu55QVaf+MUsBYsqJCjWK9eDawxOZXxudZ0HLvds9lmcWKrj2/ur46Pj05GD/d774G1/8bbz4PNu39QkcHWNm3SyvtgfGr8Wr7YRp/fTA9MD0wPTA9MD0wPTA9MAn3wMdMOdQcALKCm4r+DL4sRigSWex35JgbRGkNU2PafoQ82V/lx5bwVWBFRXEjSAtQVfJaz6O99NjXpbTda/96bHKXernNrbQlIgXbG4dvTpeur563/Y3nfWlbd3e8nRRf7ZtBNM0Lvk2D9ssy2vb0zTLum3Pnz/HwE7mQN/2dXjBj2DWrX7NNzrX1Jbu2JViQL6UbzsAiZ9Q2Je20vFmzdsDLdJQMhaQwKsyUufescv5veVsqTdefxidicfT337ucV1vfbq+9EHLifDx1W3tI6/yDNqBHwQh/Fial2Ma5Fu2SeN4S+vR903X/a33kg7JGfvdvnqMvPr+5THyb1le+77puk1sSN16vm237rV5e+02x3d781xeve86h7TjS0AjzxzjBqws4JiA5x4Vs8iQHn49Zjne++AqULkezs8uV89POXwfIO/s7CLr+OmzZ6tnz5+u7p0crX74hz8XcGzfjCVsENTqIi/19lrZgYJ2Y64harnKaXuXY71vmqyP0dm+WF67X/pl6fG9/gV7LU2XfhodfyjwlKy7ymrzGQ1fFmPTW/fT9YxHpm2tT/d1vSTWd7e9cB2LXYDUdv3hJ3xGZmvkbHSv3yV0hbzO5wOD/+Ctt9/47dXt9e+ypJ+bRQqnmuzNjC41mfevmgdmBtmrNuPT3umB6YHpgemB6YHpgemBu+KBivGIgmLQDuEj8VEiP2JQzgEiKLK6DUYN8g3yxsCXglQDYgZIknGE0y8EcwaC8vOzDMqVbsBWomts170meIyK2y/bkhk2dLEnbcjosbZ5bwnvxb3tlfFkEChB0aiXxf40qy92aVZ9pVMSirLoI7gklB3ZJmV/8a+z2douqCOn40jlls5Ksmx9UPXtt/zMCIpSBNpqpUrAEfGleVvKefrUY+Qo+CeG0ebYpJLpfwEy6mveFnm7p37OLxYSKKdIS8n5YmS1RGVTawS+6Ku/Ct6T2RbHlGwPSV/tcCi745OdUxp6xpOZZL6R0ZYAFfrZ4PzwcPXw/n1sUBclF1hQOtKm/jmrih58nYPDJaOUnLJP2+tcJoGXkXnTtkMpv7w1EhlrdLlsdAY+9tUcDX1p208mnD7f9vc85q2kg2f0QI429TpVD91Ic3hLg8eHjO29ci1ZO30fJxStftNm58eMS7XT57ccOuWZYJ1xFttp72syuEJd/CMEPrXe9VM9I233xi51QX7zqVWtHchGl/gbGoHMA5CSAsGcWmVrhXTSl1x+TzZZYtGBL3m5DrjL5/xyzZspPTfvYvX0w48AxC5Wjx8/Xp1y3tjx8fHq7XfeWP3oD3929fDBfXjpi/Kp/u7fEN8KGX76kE/WG+w7+8rn7uOy5hwfTbEZkCc+BjKqrb9wTHGdaBP+35YCwvWV4/iFil3tT5+VzhjzvtYFVyh9c628VNWVwObQrJFw1zdBianhoohk3iSVNyeAZT3oZOv6InNnXT0BD0PHb4Lz4b3K+zuurWXvWNNmjXEGmeX6Sh2Vx7OjaO/BvPTfHr8R+4f75CHyVxmDX3/3rdf/4PHjb32VHxEdz7GG5sq5Dz+qhufHfbUH1WqWu+sBn+5ZpgemB6YHpgemB6YHpgemB6YHPqke2MQtBFTGLoQ5vLeMKKkC4wqUNM7uCvYI1AU4PqZ8JxrbE8wx5uWrbLpNOj9dEoQu6t235NdjWqfvxMv2Hud90xEOtrhct+3b5h5rS4/12n7yupRvXwJ0rstS/lNeyTTQt7QNXi3Nq69p5MvAW94iN17bnubjoeYp8NkE6TY4XwTRa0EsAaeRzeJ4ZfS5YBlLfXNoP/2tm/L8oyFtKJD7jPHL/gGOJHMNuoryq085ni2lHju+WTO23K4ePXwNPlvAQzpl9Vv0Ipe6/rTY337qPtu9DzjhlSKNfmmaHm9d74d+0EkvX1ozru5t3dK13B4XPtignJrXopeuaZxn+7v+Mq0jbOtry20ejstYAUrBQ1xQ9N++ZltOyxJMSzbo4GF/f5TXdC27r80nAGjoao1IfwBq44ZF9RASM1HMw/j97FLZ8qyMI3m6BpLN5k+Lo+AjrHQJvnLJQfyCY88+OgMYe7J6/MEHqw8//BB+O6v3f+Cd1Q/90GdX9+8dBxwzc6z172vWU4TUV8+R/RbBUtdA1/vafpbGZyFrA5nOo9sjLdqkrrZxu5Ftn23y+LhfwfZBX1umV9t8RszAM/tOXx6ydbHbnWO3njb4GVmO4UZb1ENaeQlmWWpsVby3bGUVrW2wTZGH+u8KvrWftIWPoJvF/kPAa95aCYZ9uHtydKi+Tzhj7t//2q9+/su/8A//wWVRqlprMlrm5ZX2wMwge6Wnfxo/PTA9MD0wPTA9MD0wPfAJ9sAIhrDAqMraFQGTe+U2PQRNvJwtmWWbwMzuDsTqWoG3QZUBVwddBnn2GxanbXBVmFkkeTObwmjocdI32GPQatDWsiBNCc8hp2XasWz3vuvdFyMNLAfPZb80/ZbKzrSpNpQesswMckxHkYa3ZpDdkntnSR/X2CUdblWWRfuSoQFA1NkdfeZZstBCX9lV8vFjSob2rQW0qMsjuhPgdmBeB8KT3XFwFL995StfMZIuWdD3uCjBGyNveUtgtkPah25801Xz5kQIHSUbxawcgSx1DzhDVVvU6eAg7HJmGRzoAFQARBgAlp0J5MmGiZ6M0RfqIhB3c44e8gIkO+BsqQf3Tkh+ecbiQzf8SUdsXe0d8L/9DcAh9hYe8OmiT5LtFhnbLC55SGuWU9446HqDZg+evh1RtGAHgEYP+Kdt/QbSAnsE48a6VXdNEOiBR26dF+22jjrKytwoM3Pm6NLTvtBB+7H3Y/zLfcr0OTFbrBSIStgrrFIyuQSoivxoJs2Yz4BR2IZc7XROWscAZ8Of8uhiv+iX/HKmFle0z0H8bg00W8ysQ4ExzEQJyX0StvYLftnB0BRtj208P27Iwxmrq0uBKzL5Lq8BxZ6uvv71b66+9a3HOUPvjbdeX73//jurz3z6/dVr908ASh2CBegmH8fLGm2GgLpEmejX67naYxO3apnnCV7hY5v8BioUc7SXz65n+g22yd6zfdT5PSQri7XEW1ur1DpXx+gGrT3yCS9G+kyV1pnU8Nq/5fdj37VHRp7PHnla+grt88nCUgDPhWtPXsrwz7eWikv5tEDA3KqdflcF6vBbj+fW9W8bOV7pD41cGHPDSzI8a6y2FUMjcK1nQc92dtY7gNR7gGQOudhd3/y79fXl7/13/+3f/dZv/+vfKH8MnST4bmUr/btRzv5PsgfGU/lJNmHqPj0wPTA9MD0wPTA9MD0wPfAKe8DIyo+xllkBlwRiFXdRMaC0GGAZaHq1GKx18b6CNwKzRbu0/ZFWXsv+5bjm1TTNr9u9fhz9kn/TflybfbY3D68NFgwTe/iGRvoOrnvshmjBzzb7u8jb0mNapm3d532X1kVZS3/b3zy6XfAhe5kW8qTzgHOzaZ4+P7Wa4pjopT4E6JlmsmkEHvswbe+VH+1zJThvoGvY0bLDlLZeB/GfA/lEVmfDGfHbrI7jnkrqZSP62MfFLJVHD9HHw/kZIygkTY8Pj9S+3Xfd19fYAd96z0QNsi02dmoMzepqe9NT+7Z5aZ4CS94LgnVb6+a1+Xj/crHP0uOW9b7vMU3T9WW/XPSL5YX2Bf/y6//L3pv26pZc9337nulOPbGbrSYpsimJImTJQ4QAiYwEQYAgyafImwAObMN2kCBI/BGSvIjnF4EBy46BGImBIIYlxbKjWJI12ZJJmZRISqQlkTSbU3ffvtO55545v99/1XqefQ9vk5JJipRYdXufXbtqTbWq9iOtP1fV3r6rsXnl85bvoffWW163py2+Khnq6XVm3XfE3X8Cjl62CbjpS13bdrUc2xvo1jY34wmiir+cAcGf8NXSR2SO3X3rwfL6m3fYGvwwh/M/99xzy/e8+j7Ase9O5tiOG7/hV4ayldnrIzZox7jsF6M6d/uw4JE8WUo1pvQPn7S9zatv1+uifR06fg7R/BVjtE+ZoR3zkwf+qHatr+lyz7uoPvYnAkaaKTlAqM1Yyj6BvPrN0scto/rUlMGFp/tstT8w2vCbbZbm0y9dF9y09BZU68MPl2S5Xeztc74c9l0/2Hv4zO3bv/lLv/DzH//Uxz76Vn4i9EtQwfr5kLflWp/lO9MDM4PsO3Pe56inB6YHpgemB6YHpgemB/4wesD0Aa/LPrdGcMGSoGsVWPWzfee0W9wWZXBlsb/Bjt4uZJgZKG4Ee4IOXTrovbplqvu9GwT21XbJp85ul+7qs33a0/oGHFT2Qi/olOwuxzcCXTSFJ+MZdhqslh61UGj3GY1cgg4ZYdoy/hHckohBL8CNPJTYgT00DX6DfMZAU7LGEKzcHoeEfuVOfbZ55pK0AjvKMMNof/8gW9ZO3cJIZkh00Z3ME+0S89TWIddMKiUkq0RbKBmfdjqfzjuoRsW/9jtOb97LD1hdrdrAuVgYR7c2cSUrpcZRkx7uyEtm4ZizW2yfw/Rkjzkeg3HXQAXxLsUqjnuHDBuLJzfp38wNzz0vOaPNZ2jtt2Tesbno4SnEpNpHv3Tq82uC+t0vKuovtWUOJDCLJ/PMDdfkbLCcs+bMVmmdZmxdjoWku2IDLl1ncMlRa+dJ3hpTAUKpw190BQQhJfKKq2TrT2lanlmFPCxJbGzjYDCBqLPkmn/DgwyxEr1W48AfjC8ADVO7mwwmz8FCP4SxDSBKN1/gKDOPNp7wPZIuZ2YBtCEz8ylsc77DmWOngGMn+WLl66+/udx7636ArxdeeGF53/venXPHbt7iLDvnirXu74vrojO0+HGKfnWbYXeqbsfLVsVzthB7NFaeIdjYhA22pT3ZVsN3rJVsy+Vev3Rlq/osNR+pwrvdrttzbb8+8heAQ/0iy6pvINASbbVWQq+dOth+hmZRvV8D9eMEZq3pp6ydEGhvreVkm0JbfizemloF6evRxhilsajz7LLeJceNtho/7WuadNEn+CiPH1w4Z1CcUcYxheSXcVYZmZ73b+4ffOzOG29+DCse5PcojFE2tJePo3z++Y71QN6F79jRz4FPD0wPTA9MD0wPTA9MD0wP/GHwQAc47hw6I3hyT+UISit88rmuCsASqI1Aa9vXgMg2GP1azqnArYI55Vj63nWfE9gOG9ZBqzTd1/RXZbZ99l8t6RMQYZhPk2t7j7X1tD22ty7l2q6M/SugIhKG76pfIMirS8sQU/Hq56t3ZdtmkK2uLtoBZrCcAiY8PnGHrCEKDQTkcIDtAFFIzjOReLZVXbDV0tJgUsakXCP20I4IHhp1rvXRYGP4+57+pBTB3HY2DZRuW7xEvxkz8ZuwCWM4YPsWu+hQiZcCbqy3SZaK/puxD5nKMKBvH0mznr9uX9uec9fQZAZUB3HazSy2itxtE7BsQMFGadoHT8gMrQ4rP7Veaau+XSPa3O1rGWFe/VnTqddxrdfLijTV1rm+d12Cq7rEz56W9SVtjb384VKotSowVuPXlh5D31uXz1XKd1XHv4gTnGM333LMlsqHh485Z+z+8qUvvkkG2f3ljHk8uH59ed/737O887teWgRNXbce/d6yGzhv3/Tc94dE1GWfQFIDrH0vO8oPG2SKxl4vNeb+favfPXl6fM3fdO2DplmvJbe3dtH2Bp1SH+Cs9bJ1u6YE/JWbbMfN2mlJ2B5Qz62PewB50GYbbf2eNFWPv+VvgMOxRm3vOeqx+CYoU932e8VmKtBcCBT6vgCaff7ffOa3f/1nfvoff4rFwB7pS9C/CzFFF8v2x6KNmffvWA8UtPwdO/w58OmB6YHpgemB6YHpgemB6YFvNw90ME24E9Pq71dYSSgppfkPAg0mxuye713bIYmJXA2CzQTRUBg7+VxxUAVl4BwUAudklmwBgg7ADLSi1y4un+vrdUgRBRpF+tDSv+a1fvVZOou5GQr35J91YGdfZJGxJa+HWnd/7CdSj8zohHjE8wbVRYcf+Nc8G7AKLKfPJdMCAaoElTyoTxDDYnsVMl4wsXhKnnWzbzKGQReXwqA/YvcYX4Ez6uhMj+Izu8yiXYpIRg0y90jB0h63q33xy29WpwAPfaFXr+iEsfsxu11maAsAACAASURBVGgBx+orkyVPmrLLjCHZCXF22MrGXrjYoqFDdwhEPJQZFSwOMnfkz1lg0elaoX+EzQbY2posILPfLgTxoEDHD/zAB2KWZyE5R17OkVvOzvm6nsU5sc116ty4bqMvuhwWWzT5p5kZl7Klj83xVOTEbyxqwTqBiPPs+4PT7Xj4mo8kxudqypdbh3y3+Jl5JcCotGtgAzlTClnqUS4sKo3Otq30R7VM4fGp+0WOMkP8sY2hcd+CqU2XtnoJa1xRpZVV2j/KyxpkYsxw82obBD1cg/ZfBvzDJNqSEYYg33VLxgNNj8ttlfrc7DrHiXUu7LTZkC/aDl5BsNah65ThUskoUfyIzLH79x8sd968vzx4cLjcvXcX+ovlNgjpq+99z/Jdr7y0XOfMOUEs7XWrr18wNQtSH1yM9zpZlpz/5e8AaujjBYUGB0PjdyF1pO2ICkX9Hlyy3mxxPJaspRjqOpOh5i91xlu/jsrtzLH86GFevdNhwX4Tx5SVs/uQ5LjV7Xvt+V75fVAMEuO/oTsfQYCubKefLEyth0kz4xvvjl1dyt3Y6GRQ+lyx0kk/hJ4v1/Pu+5sz6Jx7jIoM2qznNxH61Y76jENgka3PZI6Vo6C99+Cttz71V/7S//hbn/jIL/MDoh8Djuk4H2aZHth4oN6uzeOsTA9MD0wPTA9MD0wPTA9MD0wPfOs9YND8uymDzsiKmMdIk7gu22sqiLLZYKqDqwqwjIu2JW08em9ae7u9Ke1rAGTd1rIrYCu+p8lq2QbzXtLbZpG+r5bdMnxuHev6iP8S+Hcw3Dzru3VL29cyWr9ypGm6vktnX+nezkfTNt/eoEn4HF/XuNb6lNV83tfj9uB9zyAze+xscxA3obg+csulJX5iHIA8Z9AJKeVQKbo2eoYvfeY/jY8edQkSWTI29Gt7xmajfAIo+sk6lx4TnMih/IAdyiiQBvgi29fKvheef144I6Xt6PH1GNuHEnVf32ObOlOU1NKq5cn+C7L7hp0CEQ1eFGlsbLmCGgVIujIGMLKaY23q0nb2s3fblGV5u3s6xx9pevw2retX+a/ydX/AL/TKe1X/hob+9knbbV/3K9t6Rs0QK3uoxtpjtl9e8Cqh9ZjjttSUgFn0IeGUtehydPvg0dEpoNgjQLHD5a1795c37ry5PH78GCBmb3nfq9+9vPKudwYcE4cU8FKX60U9bue7aqvPdY4eaxUbYs8Yt3Y0fdFVv+09zr7b1sX3xXH3+GyXX/DZYntftnfdvtbXvOu7/VfL0+hdj51B5piUYSlQs+Z0I8fGVYk8AT6Wdcu2Lgjcz5Jb72f/h4F+7jbWzgU2OJm8upZrR3zB8pMf+/hHPvbPfuaffKn+h5H8FvhnTLqSZ5keKA/MDLK5EqYHpgemB6YHpgemB6YHpge+JR7oEKmjlH7u4GokGRg+PtW+J1phPjl5TNIJ30w0DYTiFh3LNaJcgzWipQTfXy34s88AvUvT+txBWLetn20zKPbetF3v523wWkGfmUCCMAkgR8CqTLMmogPG3IkU+1lZFe5vR19YBzLNVqGsY0/H0s/6M/Jh8J6ztLDXM5LSTr/2NGiw9T864XFbo1+bS0YIevwaYb7miSxBsnMV8V+fKeVDjYeafsU+75a6V10g4Rwg7BQg4ejkWCOhiDEqzuxfIzPH1qBmZ4/pFoS4xtlfjJl7xobssCqWNtN/VKcNYQWVvBwAXJr0l7QSjfO48kxT8cCnzUlPUgb8KDJja2/vgIPujpebB9dLJ736yC8EyutYzTjLWkJ+5o92x0pCGv3aX6EY3ofbQhtzbym/FZ85kvo8czDWpvJidsAv+cvX6jMrsmTkFln8STZU+Z0ZhtnMNVW7/U19faGo6lCYxRXeoVcaQSf1XMP+2FlqsKfeL+0cmse4x3iEnYJQlH3tEwcS3YF34GS8Zjl1pliMbB3Y69cNpXf+3aK4x9lu+sJsMotvFQe0p+42R23VJvX5bUf2YKfPudb3ZijVuW3l70igzfGc8LVKt/4ekbnodso7fKnyjddfzzbIV15+aXn11fc+kTnGz0+NBbuusUbzjqNHgNavpNY4lT10MZ6sXccbnTWvoeNZT3pG3y5Zjm120zmIqltr28tbLln+i4/S6/rGb/rGjvgDyXEZf5Tj+lOOpXVknjf923b7S1bZLQ8fCy4J0PPLgBpl2r7li3J74Ff2E2X8UJUt8hSfQrP2XYsU56xoasw9v9kGTQdLjOV9KThGJuf1h3y59GNHhw8/dnF68vDa+GJvxETa/DM98KQH+tfrydb5ND0wPTA9MD0wPTA9MD0wPTA98C32gAGW/96ujCCTKKmiOmIj0o0uzwmmqK6CUAQYYHXb+q5sny0dsAukdQDbAWL3e+/zhKSxNL916a/Kbzr7u3Tbmnddl87nausAtrjXdGs5CXqxKQH3GFPr6/HLK0hjsd5BavodzgZcKf9Jpw5pW4b3bu+7NO23ts+25g3D+GP/1atj5aOjIxXmCjDlYAKIYLMJgpzzxQAApyorR/nSt87YA5iAsSVnpTg00lMELHwOP/cN+kBfnWNWtvcY5LHOvq30Z13Ad+vWraGqQKP1/Mujr9YybGufW1/3Wb9aelz2Vb0y3xqMah77GnATwGu+ja6AhTWm9RxL17Rtz/rZNp97zp3jfl7TWffq8bRd7Q/ltIymsc3SvNa34IdP5Z/ub5kuCYvtXVIHYBGWaYBWMEx7BUrULY2AmsV66wImutIG0IPok1OyFfHb4dHjbKl8HWDszp07eX+yrRJw7OXvenGTORYh44/ytbfftfab3T2O2MxgfNY+r+7znu2j3K1v5vEq/9AXEGq1fFoO2jYyW3f0Dj4xqX5uHu9dl6z7m3+wbnzYz971efNfHU/TKe9pMrvdWQTiCnnL6HXUNN71qWXdBr0ZxKfy0ePXK7/07O2bH37xpXf82u7+/iHvvYK9/BG8gtDRMst3vAdmBtl3/BKYDpgemB6YHpgemB6YHpge+NZ4YBvelv5+rsyErx29NH1jaASjnj92BojBsToVYCFZvIBA9Wy5wXYog6kOvtTawZXZPgazBncdjNnfAVr4eLb/aW3r/q7Lb3E8aTNTh+dcBtBm8FBsNaPHbBfLBTifmUTVvwVylNHBZwj5k7YBajnijvgyev44FiQrFF4zfAAQOP8oWgGcIk+X8M9xKa+Cy9Ig2KCM+AQxu6RnXOdAckFCt0W6rSogAH1m/TgGE7MiC5+XryqzSC3KMdMkhZ1QesGtUicnJ5ETP2GnGTPnntxvJo4pIfAhTBEglKfLPiKy/Q2dDs9xhJfu+EQ6M7TGeWHq47t2G5oIwtbgJcj3y4ZdyoaaZ89D8jQn6VVv5heDp6Wen3nm1nJM0ps+cM251k4BVhzinqgFJYCbEsb86ZPyA22tFvs3JXOFLMeu//1CoMozf5WhZLttHhBv8Tll6PCANb1LR/SaudWZf1S29MWVv2sfogUbi07JbXvsRpZ3VcrTumNjJNUqHBk9m/FDrerwtdroBKuILDpz7pgTSsk8NCF33alkeaybzdj65S/6bqN/D30Q9vsHCxjr8KV1jUkpe9GQDEO3pjo+17hrzAP5v/il15e33nor8/zs888sr77vu5eX3vnCwvY99vLV/JthWTI9w8/FUrq01bVRW17L/owbPdK3GdopzT5r8QxZDHDYZ90B1rrxgwM53yzvPfXNIoJcnzjvXH0WYI9TYJG3M++wbVnz3pGt3pxbNzT2rdeqNJaW5d2+yBn8m/ketNL3/EhnJpwFjcyz716tb/u8fBlSd6j887fH96rXVQ/Ts9Jat/I8769l8Gu5m3WC7L3d3cf4/ZPQ/tp73/vez53zG4MP+eYsnbzFMUUBs0wPrDzQb92qaVanB6YHpgemB6YHpgemB6YHpge+/TzQQdrGMoOqKoneyCggTmITHVGwAZSXgW4Xgy0DKUsHXmu6lu/d9qZtGT6v27re8vu+DgqtN92av2n7bl/zed8UguK1jG5vmdrZRToznNZlLct6yTJQreBU2ug2Ph2+kWYtV5rm1RdeAorXANra7qaRrzM7SpehLnNAdC7tZhscdC3TrWeCd54tdvoYtEnQbTVvFUiPcZlFdspH6DyAH7nZkui4zSZxfuQDWFKX9R6T9nV9Mzb4EFKFoFt6gQeMSdv52KLbfFkHA2DRGu0XLCyXl29tb/nyWZfP+ma8w976sl/JaV9Ja93S9zzwR8Cm5QTwFMAadIKT4QWK8e7Vpc9qanl9t39dV/ZGfjNzt61Lj8fnbleG19s9N6/3NZ30XmsbpFn7oHlah0CTpX1cvGwrpd2tpbZ7ttc6a0z61iM4zGwEmLTNjDK3BgsQ6TLPwAv4yzy7tfLB4aPl3r17uWy/eev68p53v7y8973vXm7evJ5152+JV/u9Mr+2Y9NG+9TXZV1fj8WvpErvevbqcctXY936cC3Dvn5e121btwsCtpxud+xdmrf7eh21nG4vPxdf89vX/Ot72956u08ZXe8+aWu9ls9sbxtaTtFsxzX6zRw74wJXu7a/v7f7mGP6P8r/2PBLd++8+Vt/46/9VdiydrYvhoJmmR644oGZQXbFIfNxemB6YHpgemB6YHpgemB64FvvAcKfrzCig7MnOlbBHV+wNPwzACLRp7KjCDKveQi8gA6hV1iV0wFe1w3EWr53n7ut7zJb72C3A1ufbe/SdQPcyBx92JZn28huSFBdsg1bq4Q+mU4+Dzuptb2RzTDqjk6AEZkjp0RsaH20PX3o5D/qyjQIrayUGqsZZfSVe2Kjo4kO7nVGFWrod0xme+lPQQkBqp2RRSbIpbxAENHXQaz+3CHra9iCIHCJFEGJZIbQJwBxbDqWwIAgRmzUM9STfTK8BIjmVy3VlWO8GErALOktDpQLbQ4i9sdPtglY2U970VFVm3O4t/9kMM64LBs/xNfwYafnX+nLF9/xAmAdojyfLePTiQA2OpCSdTjk1HlUdjRYgj30OQ6vLptMmdEWDgEWbaZkmyf1AAzY1JlhyhD8MYsvdfvG/NTk0qeM4Xt6QxfQyIkYxfXsyB2fZ2r1vK7trLGWPXLaJzBUNJU5JY3P63vr6Hv6Tbtj+GxopLmAbfvxzHjXag5YXpKxvkYmlTNHg5lGVtQTn9RyrrE5Emyw9AgDxjJGM+TOAoLSn3eu9Lut0g9GHI+vVr75xlvLCWvu+s2D5ZVXXl6+53vev7BtD+1+rfKUHxtVlP49Pv+KdawnQDrdY6frWRv9TRLAw6Q8xyrtYu1JjIH1nutzaUru7lgQfuEyH8Rg7TmiHeyUBgfUWH2xU/SDztrOg/pyLhjviPOe7ctZHzBESHE6jm1pj5XcHmP/3vWzJliaV13dZ7tjkiegLs/WA+QDQFqavlXnvfedyW5I+vlnyRmINeCM7+zsJLyuVjfV85t0vrcDbM8c3DzY/xK/VT9/+OD+L/zo3/pf3/xHP/4PIgNd4nltctrmn+mBtQcmQLb2xqxPD0wPTA9MD0wPTA9MD0wPfFt4IKBFwsBtAPXVDSNMIsg08CMAuzQoc69fAmZDQqKiBNJDiEFZlw7s1kFd93nvdu9dt70DRevrsqapgLeCZ7cGdV+CxITYNT7tsa1L03lfh3N5pinjg7jGUUGtdftbZ8vY2mn/NpBVV3gSaG/98VQbaFSel/IEfpJFNvxYfW1PARXSuaXNLaNK9zI2jc6cKyZ2AKhmG0N/8803A5BlTExfHwIfo9G3AGAF6AJ0uOAw/10AgDMHBL9zC8zgTPOMf5B7wRbPjAqQSPgFxemLPGoBK2hqcMwxDHYAC0ANHgM4KRv9AaaUxBZKATm3eRbw2mJLt0+OvecocmnLmkaHZpQPhj320Xh13uKH8FW/AIpFgG9DW03Rpy3q6mHapQxBHP2sM+yX10sbLZkn2tvONI4/sZO+Ls3v84Y+OmssZXPVu9+77dXXkso229TvJUikKt/h7IuG1H79rgwvx3jKXPT4wYagr/dBQE8g9RqH9ospOevSXWOdrG0RaFSf4JjZSmesUfXUWr0IAPwYAPbRIWeP3T/M8/Ub+8u73/3K8v73v7rcvrnPetMn2ts6XYOChLTj1q3HtuPVFkv7ITod8ChtY2zWHrqax77mk6Not36Wzncy75M2cZlR1zytQ3BQAyNvNOZDBtajs+yRTx+1/uoufdZL//a+1hPZg7/bvXt1nzLUF7jOgVLsiz4esx5Wv5fdZ7t+F0wfMplBNk8ji5m+bhv/Q8nDGzdufOj+vbd+9s/9+T/za//8Z//pI95aB46YQPOlUKWzTA9c8cAEyK44ZD5OD0wPTA9MD0wPTA9MD0wP/P54oMOtq9GKoIRl0z8CqK+0qgL8CrwMqurMKwPFnI+FBAOq/VVg2oGW9+gwsKLfZ+Wsy9Pa1v3WW14FbtXbQWXraPlfwUu8rMZkNI3O0kmohy3Jmhr2JWAc9pm9hOYAA7JJy0gZR2VA+bU6BRuOmwFUXw6U0jEyVnwimBDltBrY+3XGoghV6iRjZHxCWJYGixoU6nFpc+wmVE19yDoHZHjrzhvLo0cP0/788+9Ybj/znF+WCxhi9pmSd9FjdtmXv/DF5eIRh/QHR6gtZhciHRQQz9gMPOegyJ4BCKGuKmVEr8GzF/aYlbPrly9PGxwZPkOP47fUuqFOV4FkPdJ6xnEB3qTz7DWTWswUs+jT3fNrC9u4AOPSFBs4BS+ZVAEqAsxpUulzKPpM21JWa1D7peu1Yz8jDhlZMZFtdhLHkYXOucgWzTIHJ9ZXRBHPerpYOBkr41PmroZT1J8xsz48Ww0JeR4OH/6gTZ86l+FS97A3z6W/59674IT2a8oedctYAlWnTb1dyu8lPfMGr/7KGoco8ymAak2bGUO4AdAyHmSd2sZdsEsbWn7XnR9fkwKNFFK88p/jxPg748J+pJ+xVs8BZOjOGXIXrJu7b94NaAvYsrzr3e9cXn3vdy/veOGZ0sX6k1bAtuZpnDs25lbR7Pnb2JVxthtNxaS0zY4t44PeYq99vrtrwMses96cD99NKqHOWPKe+ztGXywqWY7XNaEG3xjluh23EMSyA9Zal2SXpR8aZVbmoGrK122v0roUXdM7Z9o+XogmSlvpbnq7yAGNPtsyEu/Ry3Kmf7Ne6VS3a1LZ/TtfVCbkXfBhll1+QlxHe4f47JceHT74J3/hz//Zj/zzn/uZh0l9PeNlTelJqKf5d3rgqgcmQHbVI/N5emB6YHpgemB6YHpgemB64A+SB0iAqEDPOwGx59BcGFh60HUC73FYfAKxQbseoEGkxeDaegVjFbxZ7/7maX32Na283d509llaZj9L1/XIrgj2K/jlldYgv+V77xJ9AAkJSBNAItfsmxFQdsacwfrattJtwFljbXm2N511g/GrZU2jXSWrqZSHLh4vyFr6/Gv/ZvnX//qTy+GDe8uDe/eXV199dfnBP/rHlhff+S62mJINBoB0OmwVpPkSB6G7fZFO+gyaHSt33cigYpuDA4R4/OjR8iwBv2NgTxU+Uhz0jiEPAAKAHGF2HJEBq9u6YiRgg3QBG2mnZGyxvuqbNnTKbtaKmz+19fycA78px5yFdnl5k1qBK1lvrCFt9Wr/tN8yBkRUu7KqNJ1PTbttKzmZe9cq9m/70CyARvsGOKXfzJxseaTOrOBO7Wldfa+x1JMuLoK6P7kWpFmPx+e2odsLKCOzEHCqZdW63a6T5pG/S6/tfv6K94WO8Dlvo15bDQVEmPOM3bPvCixTngCdPpCvzrSq+cB7eR9dU9UuYFZr/QzgzDn2Iwv37z3ky5UPwv/Ol18MOPbiC88vuxz8z8JJ5qIf/kBK+V3TWIuxffiZlqH/yjqwg9J+817+2o7P58x3kW7k2LYLCOt8q6ZANH97tvJkKT+XIeUDbShhpQsaHktPAVrWi6/5i96/zWO95XVb8/Vdmp7DdZvt2u8S7nbpcmC/upnK8wHS2S6tdF7FV/b5TOGW50veuX3nm9PHjvd3dz706OGDH/uv/8Kf/ae/8os/87mAYyKAnk8GZFmsss8yPfB0D0yA7Ol+ma3TA9MD0wPTA9MD0wPTA9MD32QPVPj29kq+Vv+I9wwUU73gq4fgQ6eAGNQAlUSGAERGQLUJtjoIVHMFXobNHSxWNooBmnwjCNv0r3mbp+V34Bji1R+DNwTlSB2/vOdX50q2cdsAdSrYC1fO4KHmqUEpZtPYjxy3gSWVyf4ILlk7ZFZswLHwGqwPIAWn6CDjRAtx5ygjAKWzbRfkEFCxmLlUAWz5RuBjHdAKKJhNprwGhtBCltXZcnj4ANcfL8/xlccFMOn11z63/MLP/jRf6NtZ/t0/+SJZfZxhRl3Aya2Uyn3z7ltlHPVEy9hg5pi+w8CaK8fgo4E0AJfZMpfYde6XPz2A/RjgSiRA8MtC3cf2aY41Eh1Ju75Tlv3MdcAzeASc9Ddk2qXcZJjRcCFNxNKJXs+p0sQdstXc9tnFdfUVmTTKhcCzyJTbX84sXYxPX2hLzIOWe/qGPrPHulxdh2lnnTCaVOULsOrWylXJkkHTukjbZVtfKaPTdlu81yH0pUc+fes61n6dFhnYUgBHgbttb8vve/iVwdXvYgO76UOffnIucF8IlSWthZ5l74AtjzzmXCvbfO9jR8nFIHwhgFkAVu5o1AZ+MVinlVXmXB4eHi0nx2fL48eP8xGKd73yjuX7v+/9y/PPP8taZ60BislvCQCJVypLs96ldNiH3zN/1M1y03u9BXadMdr0jqkBabdi++w/bcxWYO54IM/tJ+0oHxe9E+SIlj3/0ua/+GH0x1ZHvC2Zh2v1rrRPe27ktbQO691n3bUkjdmI69JfX+02E+aKrzULLI6xuWqyKEuGGgNs8tvgRxIs/mbmYwoDsBfYvOAkMRMKeUP3Cv8CHLvc/dDJ46Mf+1P/5X/xUx/7yIc+xQT5ArdS3B4nRub8Mz3wdh7oBfN2/bN9emB6YHpgemB6YHpgemB6YHrg284DHbwNwxLJnQKO0H7CIc2n9nfARz1ZZsZHtnexbpt063aBBcu6rXnWMVb3d1vfbe++5lvf13TdvqZv/qt03S5PgxS2AUnlalkDO9jY0LL73nTKt6391Hf77VOuQb7Fw+QDDBCsytOy9NXWzvoC4NHRIdk39wISfOAD37e8613vWn7wB3+QkHhZPvGxjy+PHt6HBx8TGCtHPcp568498TUuKNUPABBdDmg8V9DL5iwO6D47PQY0UcYWkKh9kMgodCl86ywxepzYtMdu5LYfvMcH9o9im3ZoY485NtN2esJW3hMAE2jlc0wNWkhjm5dgSde9W1qWddtapvzqfLtL+nVpOd7lsXjv9oAzjgH7LdlaOfo952t91pe6LfI2fxqe8qd12dX2N5lArWVtx1V5/Rw5w271297yut5ypdWXBwcHuW4cXF9uXC9wbO1XP0zgOJXnuhLI9e6zl2ePCar4xUqzxU4Axh4/PlkePnyUM/AExwTY3/3KS8sHvvfV5YXnby/gn6zLWutZ8/S7WMtGfV++U7422t4AknZ72Zfxwmm/pZ+9d5vtXY+c4ZNeR/laJ+yOec3ffFdl2W6bV/NY156WL43Fdsu6vdu8t10heps/0jWPJF1fy7Td53pNS6cHEep37XK7a9Pkmflr3eOO2Es/W+yYLvgfQz56eXH6D//Cn/8z/8/HPvrh33ANBij17cyY6jc9Quef6YGv4oGZQfZVnDO7pgemB6YHpgemB6YHpgemB749PdBB19q6N978slkepwRMx2bpmIAFHelkZFoYsBIjuQ3NM7oMFC0tp+8tz6BMGq+rfU1ju1fT9L0DuQ3dAFfq7B94OrgdGRLStazw5It6BqPVLp/hNJzpNlOn6MWS/CKmNhp8SyWPIEOd1cOIQ+tJPR3Ey6uNbacgSZ1NpnzrERM5YAglS7n+U4dnDHHbx4X6qW13y+IXv/CF5ejwIQEuoANfpLx169by3e9933Lr5u3lB3/oh5bX37wDEPFwefaFd4bvAv9eYOvrb3wZvsPoVxNKa86wVR0W7c0YBCPYYnl+/HjZvfkMgIeBdY0pHoIng3CcyEEA3GZSjXHjT7N1rpERJJ08ZoipM0V+SvyEb9tXl9napn+K9gLg5d69e5yp9kpo9vef/Apm+6XORlJ2yb8c86srpeni+rF0S/RjX+A57Kte/zpBBW40v7L8mqjZSZt9ZL2OIpcx05cPDbBmkvVF+4ZfvviXvnHXlir6rzLH9LNry+K45HdNeNf+nqP2WQjHH9ssAkehF8hydIyt3zf72yblpR2+ll1y1V26BKtKp87UKwWG0RgvKctsQ+n0v/IKFKysMr9WaXbZGVlj0ZsUw2W5ffv28v0f+J7luedvIccD4dlOCxiaw+EBX8zy6tnKb4u+VMNIc/MuCHfumXUhZAxmNFGcUY3Vb2X7ZsbttIc5wG7/oThj0IDIZoz8bsQP0ejyLn7XpVlqkj5Zeg23nvLxNY7l6g9VRHE0yql90hQgaCak+vSdpf7Cof35Z4blkA2dGV/aHH8qB3tib6+TsS79nGQVYTHGi/zKmnWO6nclawAXaoNbp7HhkvddE3b38ef+7h5I+eXHX375nf/oL/7F//Yf/4tf+umPezwbP0DKcKHCDXmrKoXz7/TA23qg3uu37Z4d0wPTA9MD0wPTA9MD0wPTA9MDfzA8YLBH+HRCUHXotisDNOqE80RtBExmYKwDt/WoDMQSxI3o0udNgDeCPfstfbfeNF23b922limNZU3T9jRd9/VzcWz/apcFazeNymg+G9+O1/bu9y4fYWQCWO9djD/FCYxC5emA2C2FsGyKAW7rCnAACCUQIWh09+5dsm72ltdffx35u8s7Xnpx+eP/zg8v3/fB72cb2+Em2NaGUwCKO2/dXY4esUVRG8cYVdT+cbjWU5L+w6HqZPoQNWMoEK2vzgAAIABJREFUZ80BmGi355FZzB4JOEY9PlOmc7MKvEs2BMqlr9bPGC30bq20tN74SuBDGYzTzKRHj7CBIjim6frDD0QcPjwKEHgMSNjb+3osuQ9aeX0uAMenkqEc2zMXzgdmdd32dennvvfa9Vkwqktk8tB03d73nst+/sp7rwTGf8UGaW2LTh0xytNkNm/Arbh+C4Ct+VpWy/Du2DqTSoCu+rbv9Tmbq09HxtgpW33VcQZ4075TvnXX68kJ2Io0Ack8S055l2SMPbu8/9X3LLdv3eA94zcEG/04wyXn6iUzSXAsft06Vzssm5EPEKvfV/t73NKtx7Z+tr6ev6Zb09SYt/L62btjaz2tW96msU8any2uaUs/N2/f7Wse6xafva7y+Ny03q+WbtOu5vWeZ3za/N3XsrSXd+rSr5f6GtBPAm10HdP30f293R/77d/61I//g7//935dkPAy5wJe+kOAEb1mr1ozn6cHnu6BmUH2dL/M1umB6YHpgemB6YHpgemB6YE/MB6ocFUw4pnbzx2/fve1ewRQDwi8niUADqJkEGbiS2U3FMhkAGZ7B27evUbwtbm3G57WJ79FHq+W17TNm/vIrNgZwaMhpDz8SdAqTeRkOAayQx5Bu/IEgbxLn6wM6H0+42E/GTUVDNpmUJlML2hyrhg4kiX6iBtDY/AvsKRMoIC6I9NsDQLW6KLHe1/yd4Cdun2oMntJMc8///zy8P695bOf/sJyDBD2jne8Y7nLlyxffvkVQLJ3cj7SXrazXfLFUUGs/YPd5cHjy+Wzn/vicizghd5so9RGZDJhGLANcg3rk0V2DvB0+njZBxxjY210ZyyOOzbV3QDZU4i0lZnNODszJgvCVm2np+7UoLXEh9x3sFlArOYaMEuwhK8eQrB8gYy5i4s/EVBMHcdktQmcffrTn1mef/GlZCLVGWasP5JZYgdBfGUBkeWHrX3m1mb7I/MpnaXmoOqVQYRfkG+7NH0J/Pmv16O8662OZjS1nu0arUWR7Bx9trlKb2eiudYij8wfq2UTfnJ9YkPGIOjh1OV92M5X+MZYum6eEEKwfQBbKxBDGT2Pbaf3fPEUtvaLsipzbcwz60Y7BMS0r8HbbNsb48okx4gCy29y9h0fqOSDD0fL8c7F8szBjeUAoPP27VvLs5ydFzkn0HKml0CadugTbUBbMsRiB0b3Wim78CW2mlEpj19AVRbe4o69/mTEJ/pODop+NF3TKu+/fo4e+NgyXvwIje+hFczdRZTbRZXZfqlfwojJH9vRrjEBvX0uv6tnSycgngzXld5ki2JJdA7SjKN9wH1TXNPj90pYOTxj4VwIWm14kOeU6QbmX79pv5lv9eVhfOc/6PvKOY2wMLcs84td5xiQ9PHe9f2Pn56d/OR7vvf9P/aTP/F/fxihHEWo8EtMYMCU9uHGzlmZHvgaHpgA2ddw0OyeHpgemB6YHpgemB6YHpge+Lb3gFHr8ou/8LPL937wBx6/8ur33Nm9fustvjh3+/z82i7BFzFYgjRirg73a0wGaAZRBl0Gs08r9jfdut92i4Gcde/SdaZa9zeP8u2HME0t1/i1y1pWy/Qw+w78E6QPvc3jXT7+punqOMr2CtIlEIiJHMjdbrY+VDs2DfvaFnm6XnrqOZ7EBQEvBNQADZ579oXl/rNvLc8888zyqU/+5vLcc88t3/XKu5CwA/Bwc7l+/SZZXjc2vjonoD3mU5YPHri9kkKW3wJ4BiqAbYmiVYBCr4TORL1Fesk2yzMAqYMbzy4n+IQZcCcp9AzMiD+FcRsrjzF5L7/WPFwbWYWSZm7Q1ZlnejNzxtqQLwAi4xRgADXDjt3l7v0HgXcE18xI8vyq5557YXnhhReWg+vXl89+9rPYt58veB7smWWGXdinXLfRZQPYWIP6NvMCjbZYX5f2vTIU43O3SRfZ3OV1DV7DGSXPkdT6rLHrG9uKp2U0fzw5/GSb68V7tzefImwXFFOG9bJprC95uNYl7xl74PSl89s8m/uws8fuvcaALNfBqkQX8+zXJB3z1XdEmdfQtXdQ9u1Qx7P8Kz/7HEDvWT4kYWE+PdPOw/j3AMyybdDlyJwLTp+zjgqoc+041i0w1T4sQfW3x77xjWgYQxCyItMVovZZzWVk45d1UUbPZ3S4rp8kyVw79viHvvbXWo71tqfrbX9eFedvMFwdi3zd1vXall12l7xilk57S1cZut5y6fDU4zvEzMXW/DbDYwHuC7/11nkOOGkdl4OpAVJeXJzx2/4b2P+T3/XSiz/+iY9/9Fd/9G/9zfPoubjk87gBx6IcPtWVIQqdZXrga3hgAmRfw0Gze3pgemB6YHpgemB6YHpgeuDb0wMjWCP4IcQj4PxnP/UTyy/+4i+e/PUf/btvfe8Hf+ju5fneKxd7y3WCUZIjLi6JrgyUOg7cBJIGXw1qWa/grgK0DggNOg38ukjXxb7ma/rIMCC2DI3yRw4BXxf1NgDh2U+hadlkXiinzxiS12Jb5BP32cbgAQdOE+zb3rZQSV3USBCsbY4NjoX2BMkK9YD5YWh00hTbBIcoxaM8n2pAfvUx+nj0buB/jWybd737fQG8nvvS68trr/2b5aV3vgx49Hh59tlnAY9usPXyOrL3sZntcIzxBJDsXp8/ZlqL40R2gC6nTNQrIJmq0SN4Jh0AGYjUsnP7WcbOSVHICQDD9tqLy9OFvXbJatJiRoOX8Lv+0XyWTH1FEh8KgjiwXNzwTUAynhPsJ/MnrPyBNvE2+ul3C6mu1Fdus3R76Y0bt5ZX3vPuaL1x42D50K9+eHnPe96T89iU5zzo9+jUd0kpUtxYL6wbvxiqnfFrTOMPoIL8kktq/xpQEG+jCZ4CQwUMit5WrTb0gyiFdTPk+xVGi19ztES2NsIjeWPK6sp828eVNUGbnlVWKccXgh/O07jUrdGuVAErZgkOfMwZUurWbtengNWZXyPNdJMhxXMV+fWS52txz/iZb9aIWUcNjDkHXnknoBP88lnAK3zqYYxq16Zd1pHnWNV5fTyzpsIb+YxpqPf9c/nljDf43RLc4/fuax6+yHUs1V9bduUd72QcVCOKbwTY8J5Ffh5jZ8+RsqWzZB65O6e8MtEvwJozFZ0L6KQJ4KscDfY/21uvw6ZcjK9WKl+T93i/omfoEvxaj08es7iUr4isL2r6Xf+mnSUke9usPNd4eEXgMpYaq1KyPRa7Gqyv8dUYzsjQ5H/VyEcwkJcuM4GVzTt2cXB973du7O//s73d3Z/80hc//6t/5k/9l2ef/Z1PoqrPHIuZ0c2fMep+nPfpga/ugf7V+epUs3d6YHpgemB6YHpgemB6YHpgeuDbzAMGTKNQqWDs7NGDky98/vP3PvhHfvje44vDU7LHrp8ScBGwQX4lsCXgMzC12Ge9ArUKLJt+6NjcDP4CxEBfgWDZYd2ri/wpo73ltS67NzQQdl0ZbYf8Ldd+6x5Kf0AAqari2QbSLUM+x9Pgge3NH6u0yX9Dl3dDyQTq0OoVbUg79Zbrs4CJAS7U1N1aVRlLGmTfdTKnvv+DP8C2ypeXt958fXnppZfIqHoufQbUggKX2KaEyEPOEV8gTVbWOXdL7xUDfbiWLWrOb/nWLZIBzU5POKj/aLnJJwaPRpZJMn3IKAqpDqaScStTJCN2U0e/Jdkrjn2Pi3GYubYptndR1ni+RibYpTow4/79+4PCtbQLOHZjeUwm2Ytk0AnYvfjii8uP/MiPbPzaPo0P8YAgl6X9W7aWza3P/swl41aHoELT67+akwLzpLM0oGFfAB79vfKHdL3Gmr+3S65lK6uGXoZ2X99LX717trUs75a6ayNyOBTesqaLHBVwXTLnRd/34hcEsl1d1V9rzoy9Pt/NvjqgHjpwGPW5tVH6tpXW1HfRI2iEB1TLfS/g176MtInnNPAkvyu25m340DWU5TDkAR75HtD01NJzXraXDyTssWhXF9sECy2MOvb2vXxdfNJ5bfwnPc8W29RZ213T9BV/pPFay5THZ9tb9tvdFXi1r/laWfev27uuLiwogI13Sd/xv2DwenJhQ223rLHgW3C/AuKQ+dm9a9d+jq2w/+/R/fv/6s/96f/q5DO/DTh27fIAzjN+G8p5tCiybZn36YHfrQdW/xfgd8sy6aYHpgemB6YHpgemB6YHpgemB74dPBAwgCCoYyLu1y7Onn/m+Yfn5xcPd3b2SEYoMEUggrg2eITBrMGbxYDN4vPTAsR08qfpmqYDyw74Wl7LCr1ZHKsiTdN7z9cCieE27Qam0K9pZG/Z9mm2z56xJKYDZJA26YS1irYAFG3tspGhACijH4QnGSzYmWwm2gOokQFk6cyaPEDZoIF3/BtdAj29xY1otwJuAIObN28uN2+8a3nXu75rHGAvHRljZPyom1FE58HBAZlgp8vJqVvEyAxja9vCIdsZlHReAbWw26rQhplUolNcF2TOCXSsSwA4GzikSQAsfPqeJs9Zin5AEnOfokcak/oEHVWJxGAU5Qae6WepxWdkPO1h8/nZSc5Ie3xyTAYcYtj6dUrfLtlrro3Dw6NkjAniXL9uttw5CW1kR8X/GqdqFMQX9dxrSnBQkOQaRympM2CkY4c+4CAWMVPYyNwnOyfG0a+PuBiE9a0q3xOugI3Of5UGQ3ySPrqsx5/6qegE29LHc7KheFa2V9lXdBlb5qt0bGTymLWYt694fN70Y1vkqVed0OW2AcxKfv89JjPw6OiIYRaf4El/UCFjQo62MA3Y57tQ9pghp71ZE1HjmMu2+sJkAUQCaNLhCO4192Yo6uv4QpDSLLJTQCiJsJaT42OeX8jVrhT9TQUJkVegMnXa826pY1VwK8W2kuV7tmlBfiC9MQbbAyZlvmvuCjg1g8+x1+Kt+Sk57e+As1FWc8xfdjXz/pmZqT/GWMwM7BJ/8NDy+tn+q/XWs+6ThtmSuOaasQrgJQOQMbkepGlZ3C/JGmM35UUyx3aYE5L93uBd/zA7sP+/N7/4xQ/9N3/uTz/4NOAYQ/FYR34S/U3YlK3xm6ZZmR742h4Yb+/XJpwU0wPTA9MD0wPTA9MD0wPTA9MD36YeWAdD5wTJh3x17pBIzHoyQrCbpKX6f307EDOQe0pgliCtA3jH20Gb/GsZ8q/7+zmN/FnTrnV2v/Rea/nd593A/6nFYH3wdn/rVpa2W1qud21pmid4COibzva2x7sHkz9NXvvGPulan/S5AIoCSggAEaj7FUEBhQLfUKL9AEpm/BjUHz4+yhUcQ1CADC2INEaTPJ2bPzyOyOUCPTlmiMyTk6NHywn8xM/Zlug4264wI6PnoccmZBHMLcIdA76Jrwu0sdksljVfSPGrdI4jfdj6iG2emtmgnKDV48cnyxtvvME2U84nkwc/ANaWL/FZF+30UtZal23Rx31rc83n2t/lnSfnuXnlL9BTN9Ya896ldftse/oEdIZ5V2mla1vzhdABwrWcltF36S1bOa6/7dq0Xd+s7S2OLU/LCgA21q9nvPkV1OPHp5t1J137MDaO8bRs762r25Qpn8/0wl/ac0B+xla+l8YSHSxnli3AdG3dFFTzAP3ud3wbenmGTIGhja6nzGkEjD/aI61X27zmtX+XteQB913WdLZJb2lZ1rut6/bJV8++p1uelieNl6VltS29Xtf9V+v93PzMNp7eymz99re8lq9K2i7dtizWx7y8xZx94vjo0b94dP/+h/+H//6/+0LAseV83w9+AJafw1sDUuAs0wP/lh4Yr+2/Jfdkmx6YHpgemB6YHpgemB6YHpge+KZ7wP+X9Wn/b6vx0FfERBecd3VMMHVMgCZUk6whwuEcZmPQJjBjsb4OzNZBZPfbtgraNgHj1X6fr/InK4P4Uh1P9hmMboExeS1tT+vbBJADuKhYFXsGiCGPAadFXq8UgucL0CY3G/WGI0EdQSlBKO3xkrpFhRc9LcN7ZbCUj3yWV30Bulb6BBvsBwrifCbPFDvj4P0T7qfJmjKLz0yrY1Ktzs8M8CvLKjIx4JTssaNHxxjGvHAls2oAABlrFKMZOZUlwsA03E4O6T89ehzQwq8GAisgA98a8ItmUGzvoL/b9LGgGgL5D9mCBQOUCL9jhc9iElEGzy320K4PuvDx1OXg4Hp8KoAjgHLv3oPlzp27BPaMxzwj9Q0UZjMGvUlML5DV51aVT1wbzt8F52xpu+F/zU3WhFljYobwKdfLeemSudiAH613+/40ONT03uXpcZcNyDZDK1layhYcrC270alGMnbcFqnfpBAcpCHjzBpzjWcBjnmAKuPFNv3HyxmeHv/GDirya2dtm3R9XeMcOwBRruMjtlayxuTTloAo6EI7Q2C81sZazriwVfv9LThzrvU3NjiXXhkC9HsAXjEK6ozRPuUis8YM0MnBZIKdzrHnxFm2/mTszHWffRYehu49clyPrk19TXHra6qYdzHOz9Mu65fMt2suc6Gtod9ugbRdHyk7azPvCDzKlHboyFip2xZa7s2nVfbrl7w5Dl9FK3/ZFxtW8pQTuYNemuLDFOi6v/kig3Hr+9AO+qxltO3hT8X3FtkII43NIfmVzt29g0cH+zc+g+8/TGbqR370b//NL33yEx8VNPPK0BAZ3Vo/y/TA1+OBucXy6/He5J0emB6YHpgemB6YHpgemB74dvCAQVKVyiI4JvI9JhAkIiO4HAFdk7itp4NF27puQHe1rNsSVBuQUuRpPgPOBLYGsrR34GegLL9gQAelzbuW23IimD9rPd0mvTK8a2bfbeMpZC1nLdsOn9uuoqnnbJdLX9gZFHcutyHCED5t6a1eg2ojy+eWXT4oO+ILO4c/dgRS1EP33t4BIJoHsZs9poAdgDO2WJoVBugQEC/gQNmgvSXV7gL1lMMGLOQDULCF8RIw7hpgnEDJGbwZo+OAPl8LFJhwTJbYBIDoGWKOl8A9OtBj38IXD3MH/NgZwJ/+RqHcgBdnACCeAwbQh77jB8fLYwCymwImAK+O3bGaWeY622c7pmex+QXE9lVt+6v5jEx4Mo9Dh3Tr0uvBduvCNhbnqfXl2TFcKfL4pdBkOgkaItr16Jgz7o3MLWO3b+0te/KsjFWiTkBGxSKntjVu16MSsy7oU2bb2vLXZ6N1W1shX18B0xi34GP8enJeoNigkUd+L8va7gKvAMZcX/gtfg4A5DRX5ljz1nOt+whCXsaFHm0QiFrrQAJkbg9M15Bd+uV3/SEgV8CoMi8ybd7IEtSKj8omaS1pq2qeHV6PzXHUmMrHthdRrQnH3W2xo3oD5snXfQ3CacumDdon62Vrt+mn+AydAmNZA/D0eOxfl5bdW3UFyQJM6h/KBe+s43GLMrSX2B5P6W7q51z3OVvwt3hfP/Sl1z7/iZ/4sX/wkJcecDVwmz8Ea3WzPj3wdXlgAmRfl/sm8/TA9MD0wPTA9MD0wPTA9MDvnwc6WnwiIBqR4bCCKA5gwq2Vnklz0WdODZCKY7+MvbaBbtveQV0HeQZstnVQ2EGe9Gr3uQGmBM+jzX6L/XCrimyTyjS56HSuIkmQiAIizApONU19bYOgTuoVL8JVQzUbpT2R/uZLsI516Ivdg99MC3kZdf4JRKUY6FYtAapfxTOTyrFbzCoxqG29GQxPbV/7ps5S27Z7UP4F256AkMKqvzzXyfHYzhP2kYWlfei7e/f+8pisoNgFYGYJGGYATn8VbMNB6jbfRbAjM8EZZKdss3z2HS8vFwBUZxfHka0v9SufzCRFDdn6eZT4OGNUFgXAx9yffDjAOTLriw6zePSFJsmTTDLmQvzOr+wJzmnP8TFjuU6eGNlFAmhmrwlCHPMBgdOzFwHQHgVsi+3Ob7Sh16kaY7pqX8xyrNotcBB7K2PoIoCjfqn1GR+h07vyXJd4OHOt21tHZNFnyXhSY7jI7rXe93ThF9jDH97oo6EzpwZfyw9wFvE1TzCWGByWbLyMBbDKZ8w3K6yuACPxkbbsHZCFhX8FIi1mzx0ePloePnxY4J4ZXOOst9atfYKW9Vxgndr73cTo8qUCyywqniFW70p8SPslkz1WBf0lz7Wq+2tlItt1i79POSPOpejYsk5YNNEv5airLr7WtqHYrLzyJ2SQXrjY0IVYnU2f82pVjppz5VjyOgr6r8C66okE/mQQyOILrn58AMNdD5bYqGCKsnNeWvRVW7f3vW30OfUYiBzlycKlT2J+Efk3/dJ3xqEqS9bQA78Zbm1Xf3TC7FJBUxE3NFy7vnsg38X+we59mj57cPP6Jz/0uc99jpcKB11wBGOc7LTPMj3wDfNAveffMHFT0PTA9MD0wPTA9MD0wPTA9MD0wLfUA26lJKbON/MSOhkkGxBaDIQTHBJVVdBWtna/bR1IWv9qtMVZf+WxXOVpfvsSrA46ny2t13rzXq0neB+0Td93ebwstqmj72aR9HP3h/AptN1fNhbVHiCAblNe61jTWY/NqF/b2DTdbx8hrZFzZNlum/YJJj3kQPtjDgknJSsglQCVI9ojQ8ui/gB1Y5xmdqGZ/xBKJtgFmUUXbOEEnZI4mVzye9C940kRkbE4oJXP0kZQnnHYZ4FPnakO2mzBpEGgKv7AbssZ20PdTtl+fuWVV3I4/w//8J9YPvCBDywvPPc89FgD2JRxwCMEY8mzhq5K2xEdY7z6ydJ93nPFBsa1yuha03W96X1OGSDk5nHIU+fGX3TGPtrkt3S/z9YtPW7rTd99tjXvum5brxfr60t5Xlkb9PnuHrOH1eyxHOjOs5l69vel7La7ZSt/Lde6JXMx7hkPgKdLpG0ufu2ucStn3ddytKvryi2+lU6nZfjOu7Z67yt+G0uzxyxgVF4tecpUz9WxKKMBuMjxeVViiwlvY8zewzPslHTdt2JNu7Td/wQtasTfLIy0KuNvt3u3L3d8p30ta3233s+tT1oKgncuzTS1nbk+xXP3+N86vvSZz/zOl//+//n3mBBItGU599PET9gxH6YHvl4PzAyyr9eDk396YHpgemB6YHpgemB6YHrg28kDAmQXBKQkKdRB3iMY42YCmUGoZ94UsDD6NoGrAzEgtVTcSR4Uwe0TdIRmCeogMBPCrZTyRDZtTSsQ4hlMZlIkY4Lnpmsa9WxDPHltGcF1VQtQEcQZAJNZJRVUwxuGirTBBYcNFXzuoLf0lLyWO2LcDFCbVVrnIW16Ahooz2ywzswRJJLiOsCV4xBAE7TQW2YqqUt50ruFkug1I7A9dPRpt3jPCIbDc4cMsrNzJCNP8OviTJsAn9wWR9ulaTPKslnwyryVATigcQE9WXYAyvyyJsk+yfDKFx8BjpK1J6/BNzRQp+7B3gTYwweMp8TH3h2BueisdRAfDz85n7tmpSUTDnLaD9lOeX5+K2N57rln2C7qGVuXywsvvBAwR+coo+c+SsafrKN1XVsp67WkzaFDl3I860tZzpntKdapbLJy0G/iom7dbxpXkvz8iw9LFTLlG9tDM8dX1nvbVABGqcM1giDqdx1Y2mbxi84y8ouNyRBSJwb1F0+zfszCG3yp8Md14dlevjun8PrBg0eHj5eTYz4AwZh8F/3y6fXrdeZb8RUwZV3/+BVH123mjbZdDRrFTMH2mbJ4efFTnfeWhax3kOHZ+9oirXNpaXDNTEa/mpmzwqDlO4vMBe/eOe85gJbvu3w5g5A7VpUt6PMdGu6iuYBP+50XfbIuzlHmmz5L2913tz43T9rMTHMdbDJOyx/2tZzmXbe1zm7zWC/nz+2T8mUE3AMaajzvYM74c26xHVfFdfpdHuVs7KJPPtv4L6Xl6dZNGxWs5305WI6OHwOQLdcOCiDn6LKL+5R7f/kv/U/Hv/qhX0CGWahllpqHWLhnmR74+j0wAbKv34dTwvTA9MD0wPTA9MD0wPTA9MC3jweI6dgc574oYSmDPQJd75YngjeCMtttszSNdXkM8rqv7/ZZ9xL06tL9axnd13K8t9zu8y5v80XuCJRbZiJqgtGmMSJsWRsa5DSQZ5bTOsOl5csvnxk4V/WWjzqQxnWU9pvglzJslV/Z6ccQZSmXPa30bW2URn4vSx2kvrWbjvCeEjzfvXtvyETGiHtjs9OC3ioYobsDNjZwhWxAUA/qPxcku3G77BEoM4iHXP0X2gCA0UWQAoJkg0njmK4xjtx3uTu+Mjss7eP2//npGdtmBYYAfOCVvvvUJ7ji8hPIic8FYynKycUYpbOvr/ZT09jedb8a6XOXbs8YV+1qkS5g5QBpBFGktwS4YnwCPY61i/1th22tq+8BG5G7fd7K1O4hfmvvENz03tUnuOi66PVje9sWvzEHAa3gFxz1QP6jI7ILySDzWdobN27Er+2voSq22V/yBA+32YP6QF0tmxmHjkkawFnb0XYq89ytlqA9+irn4sFvKdonf0+6XfDP4hZKizZKv/ZRt7f/e/woCrCnb7rNs7nkR2LuzbOD7aGhz3vTF23P35an9I81MOivzoG8ze9h+tGRdxFvjVewLBnP0ttO4wYU85H2vHn01Vbr4evRx+0r7K254kxCski1oj5+oP2+Jzmn/8G9O289+NUP/wqLQB/7/rKYvFNqZlKdf6YHvm4PTIDs63bhFDA9MD0wPTA9MD0wPTA9MD3w++mBEa+9bWBE8AcmwklBFmAdA7BNcJmAviV8ZbBmMGmRs87fqrpt9tleAevAUAg4lW2Qal/xVdCaAFLq0ee5RQXbKK3aldln8GzlV+DbskIs0DEC1sT2BrqYkuBYRITSdji6PbJVCKPTph0bG9qWcZdPenWhIra0HQ5VvsrAyUN80EG8X8q0SKcuBQhkyF+29FY52wx2sVlfBaTxeY/MoNPlkDPEUsgw2mWb5blnqBn8xq/0mBFjRhDPSRHzbCqvROYoNxvs/CS6z5i+BhZyjplglwaui7E1Ml0bpMIgusZBihLt+J7n0m93rYdmz9gALupLg4zFf84Fl2DhyeMCSeRm0IwUAAAgAElEQVTiQ3xp18PxL3J7jny26ELP2vLZPkGclme/dfvMDLKkHqiy+uTxsjfzpgyymwR2SkXpdD24nqXFstBuZCu/iFWxKb0OpEdz+O3s7CF5AoLQp93SWzaAEkZFrsApPq8vq+KzASDZpw391cfm7zEJjplB5pcMlXlzb3/hK4YBWws0LjBJ0+MzdSOPv7n31KUvc9FgeQFMttcYmXeK9kGh0eVT5wtZgqHamm3CPvPtj+btd8H+vswmU25cjYQTgDP9s4cfbD/jHpv0KXprZstX0ilH4NX3PB/6iHWMSvuYigsi+IB++DR2MN+xw/7Y4XwBaLMUd/b9oi22IS9f6aRdfb4bAYKV7fjKWJ9io/dkjMW3bWHZqMXq7fH681PnqNHDgHrHLwdAKiaArXe9XHz6h/dXADDrutalr3O+cru7T5Je6cQGs4GP4DvybEkco6ivXlZOXVW/Os/snR4YHqhfsemO6YHpgemB6YHpgemB6YHpgemBPxQeIMzlS5YJT/n/dA3ILAamnTllYNft9q3r9lmapu/SWO/+q8/y2Nay1Nel+Zq3n+0XDGi+7kcSeorbPrcsbvu27ZHD8NbyWn9RbW1qHd0vj/W1XOsG5DkLiT6HIPDlcy4C4wZCwk+/976AYNKv7pYtYGa/AbyXpekhAtTykP67NMokWMiAhu8EdEKLj7xLvyk85+MDIgYc1H/y6BDbC/DQ9wEaRtAvGJACv3Kucbw3FaN6LF7NK3RmfoXGngZ9pB1XvmLZQJNAGmPaM2UMNMLxOZ9uJ429G2PLHz72uuh5WN+1uZ+lbR+uZTW/bd0uXdM2ONX9TaO8bCsecut5K6OfvXeRt+Wqt2X64QvbK9OnxtR08jadd/3R8+5aiI+cbHxnkY8/8UuPzWk7Ahg7BjyV33bf3Vu3biV7LIz8aXpleCVLEdqmbzrvyQRT16b02Apka/u3trsuam3k8PjBZ3+2HIMKKVNdfW1EU+m14PbM8LA2HP8JH3bw7tW+8S5NfAEv3tnI7DZlC6SveexrH3j3uS/prWc8yK96jekqbfRD793iTchV3jxTLwh2JXP0hWD8ad3re/jH+Kz3OGPXSoa6/S2w6Dvn3jvX6cnp6cPrt288vH37tgsiNPwp4/rpyant1nmfHvg9e2BmkP2eXTYZpgemB6YHpgemB6YHpgemB76VHngyMtKSkUJFGGdcR6iYr1gSqHFcE9Qjk8GA1+BNIKIK2RUGXLB3oGl/F4M42706eFw/dwApfffLL014G3wJBrACMYYOaaSXV5sMxC1YuLIZG6CRTvqt7dpdeoa48PonutMHcIPuHca3ts/wN3RmoKQmWcn3YPsu9vmlOwSmyTB5Bx/uk81jFpEBrH3+i9/gpQce/uJ3Xa8tYl5KcAum2Tg7fn/O8aLzEdsjH9y7H/lmxUAA8QG0J/Aa2CsrlmQsjCa0CvSMNWWQCrOcHR0vFwTVy436cl+PV93RjgzPSMKq2hobmfQAYMTQkrr5W3Mz5tWMLGxPlo1jl1fdDH/v1s2FwD3jfAL0QJLAmX7xjC7tiR/whyCWvrkIQMcdUC7gGCtXvQ0eaYz8yRyivpmZ0BWoIk2KO4qTmVX8rnX90yVyM2al1FzHN/onWTxSbte5T7EXjynHLCSsthmb0KEnWWMRuWmvfnVlvJgkQGRmlr4pXnXDrTz4vXbJ5suHFxB2OoCjY7ax6ge/VunABb/2rx9seOR3LpW1GWZAK0dR73feQ1ZIQN/YWuPWpyYw1TjKZm3zPTNzy6+ralNtNdQ9rvuam6xzNAuS+btSdJ6dVXN9yrbQnENGFqQ+kF7g2LPwzCjMPMQTyMWm6I0PPJ+sfAJZ8eI3/5lAaRZdxoxPcnf8EGYsyofXdeW8+I5Ks5l9ns14JIUMyjifOwX+vMPWKb63/Zw1pwyVj/WhPEE6dSKSd0cRrI3V72vE9++L9vv++vMMj35xTlwPeT+V4zhiUq0Z2/kdhI2MPX4PeS+Od/d3Hty5c+fh4eE9F7mWaq5lU7HmmLYN6f+K52qdf6cH3t4DEyB7e9/MnumB6YHpgemB6YHpgemB6YE/eB4QATglhj8lGCMmJcAEjEmwWmFhBWcQ2VcXgRVRmnVLB7Z5WD13fweRCfYEPozwRpFm8zzktewEhdAZ9HabbFs5JSR6BDtG4Nky3Yrn9q185TGBZQXUBt47BvEj4FZK5I+7wE7b3n3pR4ft2iWvdWPZzhbJMW4wJMhFnzTJsCI/zxLgDkDrhK2JkW+QKr8+wZWeKRSbyq3h8ZQhwaZglAT7ZgodHh4msgVCgJ+A2XFI4J4rg239G1+OuwE7vrnwoPzYgtTjowAl2pJDwJCNENiM4gl5rpGRohz1I6u2lKFDusi2yz7blL8CRKTHv5b6iED5Sz/tY+fN6zcI/o/S79h3/YgBWWTq8coB7t7HHOnDa2wvDfaA2D5Tar2NUmGxU5tj9/bZuetivZ+bvrtLf1N6d62iL/O4Xe9IGDJ6XaqSfnyTuaQenrG9Tc+2rtJhy+BhnF2HKnJaRt9Fp5TdvMq2br/X4RFnygGm9Nhu4F+3VgZAXemxv3gLOBbAVQ7DoeBYFqO+rYayxZ4Cx9SvD2zpvrJJegEnwSGBRp/jD4jLptLj+netCJJRgYetxNTZKBw+abWjs8h4SKn2mgftLZnow44UX31lw547jd573obRRTv+Vt8A2gNcoxkRu8xZAcyIiz3oVfYord9HfR89226YfKj3vs2TVllukyweW8rG1lFyS6a2SZf7sCHbdAVPaTdzzKxLMTzrZNldkDHIa6T8szt8cuWLvDN3eM9OHz1+UDYFsUYnejPd6s8/Pd4tWjXL9MDvzQMTIPu9+WtSTw9MD0wPTA9MD0wPTA9MD3ybeKDjOAPjVQFf2REcO+V8pIs9AI9TM2AuTi/3ibArgKuAPEAFwWKfGWRfBYjj/0UGhPG5i18PTEmmjsGfgbNtHWBbNbotvgRqdBu4dVGe2Th1zlW1NoBl4G7AaAAcW5rPYH1lp6NNhtAQKp5TQezWDwlQPfUH1XYnQB1jEcSKTQMgEI8yrFS1BQurMrJmsDat0ljInwFgqjEJKHWGWgfAuSNsk+02hl9DM/uGYNkMG3z1+Li20iX7SVsFqLx2DtB0FD+gIHrHQKjjX7+Sqf8dk93jgHS/bnjK+M7OyCYb8+n43QqZDBtoLznKqIp314LZO4yNbKUAYYxthy19xvJZL8nsgw5H13pgKyWZToJ5jvHWDbKcTh/q5IAAyt71gH5EOvTWts/ZaykDfLPu0PoQfMG3rA8GmvlHgKCarrZdLE/sIxVusU0hFHFTdhbHnsw9IFwy1FZzrjGR71gpkG9kKMvxOh52tZV+wMddwUVsyJno8iAPS2jjPwXwLK9z7lVyyn6zpnxWneu1z95yuiyVwaXP6kMP0gYo0beOl3/7zMltwLGc7zay0BooKykKYv64bQAm7dJK5Ol/M+C0rfziHNY8Cvxa1GsfCzPP63GkoRYe/kIOdKeI3/U3xU50+TGGLaDn++08OVHKw1/wOMe+g3m/zWrDz2bVVV+B+I7R3yKg02pnwuNP7FUfZuZZGfK1nbtDtuM36029ZnD6u2jeHm8KtMikxdnLWH2H6FNofhvG3NlUQDKWZ52qS4lma5Z/pGlfa4PvY81z2dVj0l7r9lmShQi9vvFDF8l6o//o6JC2y+W4jhjbPccvJyePl2dv3T7au7735bOTk9dOjh6/gVbSSnUKY3Qw/N1aFCuiZ/MnA+RpTbTpnJXpgad7YAJkT/fLbJ0emB6YHpgemB6YHpgemB74g+EBw59VCJTD+UFHdogNr10aiJ5y7k8Fcmu6bfBmXwWNTw64AztbO9Bb03WgKp3tTaM5azrrFTCXHOWteVr+VXkduNpvaZnNa79FgMHwsPWv7yHgjzw6qWXYbluXqnfwXJFld8vj1rMeV/Pp22FC5GpP62m5tGyC8gY2lGc731JY7j18UHbQpnyj9mscxn55dsLABGeYyitFkELL4689xiUYQVB9znbN5eAmeAkAm0VEqUFNtpdtP3xHUB8QBRr94iAAJ6zHBNZDtskBaGWstCdzjAwh57H869dAAQdRdfsW4MUdASnPW3M+CijSBEEFZRRPAUn9bNvVkj4bAQHs9xIAdbyxZTAIYuRQeYAnP0rQsqTRBreyNn/E2ViQyIbWdmnaHkl6TbU8abo0bdOPd2qjp3QX4CKtYE++8ol/22+2r98311AMRongmF+u7O2Y1/evLwKee6wH25RvEWwTyAwvaJQfCqh5s29kM0JnxqWlx9J2Y0L9HpS4Tb/y/IiE0FZvNS6eiMmfrQ3t88qOst1MMpfS/r5fCm1f2lbAWPtPY9sffZdfutiAXfpo7V/7C5RC3lhTWf/6mWdle8UXLBj7HF7eFXjl9yobKrOzn22zrJ+tt3y7i2+rp/qKx/FYtN13QOArc0Nb8w1XZ9zyMrZLQOxL5vzi8ePHlySOXTx6fCzadgl4Bla4Q3apCPnB69B+DnveiMwg6FHYCKSqZ5ke+IZ5YAJk3zBXTkHTA9MD0wPTA9MD0wPTA9MD3xwPFBB0VXYHXU+0G+uZZOB/RHYGepZrACXXshXKJ9tGOzRmM0knUJLsLsCTChora8M4u+SUvA4cwwOfgWzRV2BrtojPnSESTWRjJVgVzNjY0UH0lSDeLVoEmQbEpkgkYY1x1RlF2Iv1ewmgyy5OWnNQjKgCWMdgkW5tl/pju9kk+mYE0SE2CE7F7JfBl3BVuQS0+uCCANhtdvLznEAdA83IEbBQbckt/WaKdRHQ8Rwn+/WX2TKnRMVf+vIbBb6RIWNxLgTFQDYBygCoTjBG0IM+5lQF6KWCvF22YGEUY+J2/Gg5uvfW8sytZxYOoIuOc+wyYA/z0HsxMs10aoCnkZDCxCMEXQcDFAN0yVgYfb64p+rYgN9w0C5bS89PTpcPfuD7lutEVA8BcCyex+Q2MdeG62AvX+wESFM80Eu2kA5wLl/Z1GkUzCv5DLK+Glpr0g8KVKYiY4kDQp4/6nA+q7g2h179MbKj7EvmD7Tt/7wfPqMx63r41/FpZcatXS6+8Zwu/tjXFx5ElL6udezmQtnMZtMul4q+sO5acesht+gVvPKriuoUkvL8vfv3H/LBhnsByjzX7dYLNwP4PD45Tn/eN2gFgTyT7Iy5NIvwBhlcgic5D0xgVTUYEuiI+wascTQaOEplf/pQmX94I2PhkfvwBvTyJBsPe6038OacWtYgaH4L5HENulbNSst6LFrXhBloyaaCTnrX3gVbg/XD5S5/d/3wA3lkZqzR73lg+tx5c5WY1Rf/wlEe1Ldlr3Q5L41HacywzG+auuTmWRCQgfCfYGLZkHElSy2r1GlSFQXZve7gla5t6S3Bva7yOyQjcyEd/8GOEOwe1tHmKF0XZ9cePHx0+ehRXWyrPD85O3VLPNjY7s7ePtm/O8sdfoE/f31v/8t+EOLRA7I0+0C+GIigr1Z+NzRfjX/2fUd6YAJk35HTPgc9PTA9MD0wPTA9MD0wPfCHxgMVexnJVfF5l+DQ/z9XmKOCwoAShIOJ2ipQNPjsZ4NJi21dTzCZoLD6bLetgr8KnPvZu6XleX9aW4zMnrkCM+SRbq3TkYSXe+SM8LJl2me9tyi13g7qfX5aaX77rta7LXyOxWv4ynrTxz8bV+uXGqc2FRsBvNvPEoTXOOQ1OG8Z0p4BHFwS6N8l6NUd7Xf9k4wugAQhDmcQ9CAazQxTRuxChluxcri74NY1MlfYquVWy5296yVPACDzWWAX22xRBCl/estgbOp1gDpBIUGXfCyARwRhT821egVbOiuKDbvL8y88C5ih0UUT+9CQO7rEB3Y1ObCAZNqq4Kr3XPaz2/wuB8Aj4CMeUKsvLPGDMpx7fZzswWTtuDYRzZ+WWbYgDK5ssRt9SgqN4xx1M5kqM2s7n/Y6L12UVzK7ZXtved3vvde04Jj9Fu9X6+p9/Phoee21z7Pd7gj3CHYJ4gKKPHq8HJMBCpCy3L93LzJcGZegcN7FVW+QYfbMM7eWV199dXnm9i22GZ6xzVbfMHYB0NT9Jdj6PII2z9Xe71OPeWP/AB59btubf323zzkTYNZttcVVE2rs8mf9QOD2xWyfpa3XorL0mx8Z8H4piMjianv6rDrp1OUW0vLt4BNA838I0A4X+nbq0nbVduWqRxzUubbesr3HFmjSv+lDhQgXjb4XmScelSUY7f2MMVm0okA9x4JtoOQAY2SL+ZXK42v3Hz7Y4b7ziDMIaT9o/ecu2Yv9L1wcHPzyyfn5v7z57O6XP/yhf4E+QeiBLqtglumBb4IHJkD2TXDqFDk9MD0wPTA9MD0wPTA9MD3wLfMAmAEpJTu7Blw7BqUCLoRnAccqP8IIjBiMQDr38wpgrRukGfR1cJw2gk7b5U0QTeDX/QadfXUg3JlBHfCFdxNgDrCJ7XkIUXwwoNCS1eSdo9PSjuB6JhDNoeYj2Bc4KNlmYzmWAiAgj12OJjYl8K2+klvyred52K6yklf37u/x0FnggiCPwr3BG6/SYFaUQXQFyWSIGEFjq5k+kasd8Mnj86kZWAec5UTj4eNjOvCncrs4JrO5OsLXTvtISfJeX9a0gSeybIQJQLSonwFGkcGFvwz1zfSKfvgTqMtsHzYYZycjy2eD9wTzhSik3/QnwTmKYEbGy3xl3h1vbLpYbnJGlux5ps2pE0CLLxhDppjxjBGEjnyp3FGMLSU/erS6lmb6Y4cd0NXAWcswKNuibH25ocNf2qfnPBdLgEKwr4A2wZ0K/baQm17SJSWz1rS+0x+lchi40eE49Z1rXIDQeeI1i72+T8rwfDrvgjdn+LGBpwwDftv8sqfa1X3J+/fm628ud954a3n48CFHwd1Y3vnSS8v9B4cLXy9cPv3pTy+PHh4up3yI4Qb+9tonfev5mwfLFz7z6eXenS8vjwFZbpM9+Ef+6B9b/qP//D9brj//PBmImZjocTyuG5Za/Knf9WOyRoP4SFFZXw00C05aau4At5xzmlyF8YNC7KdRIMtz6SyuR9eMXwpRloCQusyC0i8HAHoCkvEwvAGE8lRrU8DM7cd72M8mxPwe7bptk7ZkpW1GhMWaoB3IyTpwyC4PmvZAWnPeX9Y3bZSc29d2j3fB+an1WjSZQ6vQWVdWxktFVvUEGNupDDReuYwnbyx2FG2tTV/NgHzwHV+cXTvFF6cn55ePDh9fOzx8kPl2OzNA2XJAtiXbLZcbN27cfe7F27/Chxl+/NrF+c//5b/8P9/9qX/8Ezj+HNHXTEatiSlz59/pgW+oByZA9g115xQ2PTA9MD0wPTA9MD0wPTA98C32AIkVl9exwVPeiScFkepgaLfFGYx3fJngDyKBBIO+DuwSaNLufV3vsMzgVpmW5snD+PMEz2iTrvWZGWIeROLY6Cg5BqqW1qsOL3EIi/wGppbWaxuiUxqIaF0G9nBnuJs2iJ9mn20t07vPbW/r63afQ9+Bt0G54xv+ipw8F6ATPqzIXWDEKeAi3l/eun8v7QEVE7ADAghQnuMdgbJdDsAnKywgp3YFnaNPByKk7fZQcqLr5YxzyHav306fGWcCAr2tMjoCTMRd+ZPzymBlpqtRQAC9qs7WNG1hm2DGNMbNA74hW4bo/+atGwAAstZYrWX7H2BJpsUx8SXN4h+AYWZ+a7s8GQd36bAgz8Fy8GnW78iCMmvoxG2i+LFklt1tHxKgH2sEWoEa10BGOGSZUSW9cnuOt/xtY9nS/kVAih8qSDYaagVtHXdwMvwmrcX3w0vcqdvW960u+69la+VvfOJfk0H2WtY3AMnyO7/9meXho8PljTfYgousGwfXA37ueWg//n75heeXN1/7zPLojdeWm4BIN3ZPOcTqreXjv/xzy+G9Ly//wX/yny7v+/4PLufXDpYzsrq6xJf56ELZpi1anTsVdVl8FoxyC6LrtO23bwNK+UDpvn43Bbj8sqznwLmM97m73llQGV/Tq0P/mxnmXaAJzZDV/Dw+rbMT5eUbI7wLlU2Wj01ISZOyIttnGkr2drw5k4zHbctq3PAK3QpON1/ua+LI7QbvpUM/BSClZQNuD3sEBSsbsT5CsNlqrq10nJ4dg/UB7Z6dPeS69+jR4YOL07MHgICHp0ePHl7fvfalL3/xtV989ODOz/31v/FXvvipX/uwepl1ofjgv9xmmR745nhgAmTfHL9OqdMD0wPTA9MD0wPTA9MD0wO/fx6oyK30mTW2RyC2T+CYJJAGATznyMCttwDujIyaBKkDLKhAueKvChpLaAJCaAw1OxCVdn3xkEAzYRyUG/4KDKsvPNohoGBQ20GnQfUYALcNMCZvNefcMUm016wM5cdeAuPYEShEGyrIR0MFxkOAdhvgls7WXXaqb21vssfGeIb6ZAZpc/Cd0SiPAX1ZOfxBn2eVxTbtx2h68o9G/sOPpBM5H8ePT8oegSwJnQcRCX0tAOOAR2GDVoFnPo+spdisD/uKgbIjJ+lCgEnaYLu6BRjNeqJZ0Zsx49MADkNX1gSZPuvsqtDbL6iB/F0m7KWX3uFjARwBBgY4hS7Pn3IYmRufBcvijxqUgIrPOXOsmnhGtvMIY8+jYKCucO3WMGudDVNzqzUM3OEYJVpNkjoELQS3AjAORkG+tidzqP9N89qskTGHZrzJX8snd7yrldBCw79IZnxmDzrOrIi4HJCIXotmaYdflfQQdu10HX/mM59Zfv3XP748YpulZ4/Z/vqbd0offAJmfMmQ+/7y3O3ryw+8+p7l4eufX5bDu8t7n7+53Nzjwwxsn/VjHFlDAGSf+Pl/upw+uLe8/4/+8eXGc88nm2u55ldKtZRzyii4Orp2AGH1X9xGuwBYMrWSyem49bdbB+3z/aEinZNL6YxOx+1vyqVnlQVog9b59x/CJVdP5PBQbcqt99W5t6j/ZGSjOfFmgWWt7F8GfHXLrrx61XsBlXKqx7s9/q17n5nm2N2snH+ON+NSBrSuEfj9DcrvBM92bHh43mMw6qMxd8ft1yelkTY6qdcXbocNPPtlTX3luATkuJ9xft8XWCyf4P6r73nlXb/5hc99+nP/24/+7Xuf/Nivm0p2spyc3sGJb7oIMlZ+FLijSrnlpyicf6YHvsEemADZN9ihU9z0wPTA9MD0wPTA9MD0wPTAt9YDBFGiFEavFbVZMdizkUCtgqwKCq2nb9wheeK5aTsYbnrpum3Nb90A0pI696sy7Ks2bQJ8wNR+tu9qUU7JGsEoBBXQVwCLtLDUX6pj1K3f+xbgEwgofT0W+623TJ/bT7Y3nUqkCVqjmsFn8K78MWzJ0tcZbW1XAECINM++Ew6592wpdZ3aLmCkP5CrjWbhUKkrAI2hC4E69J5zpF10Kowbdb6CeEoGGegoVDzDG50JzpGHzoBO8tEWQCy8yBAsOD9ddvgKpqCYvCV/u2b6IwmG52XjlkZsqUtsGw8BEJLB5DqrjED3iFniSyuqp63Xk939XH4da1RaSuu23jZu6zWPDI++Asyo2Z0ivfwMcvuMAdkm6Z1/G/mQZE0obAAVtLBaXUMOeNwBeOLvvHKk+ACI6FZ5Yx+k6/Ukb7a1ArA41s+/9sXl8PBRZIoRCfh4NxPPtSUwY+LQdUC1Zw92lxt8oPaNt768vPMmcwgNx/Uvt27cXk4e++EHN7BCDXj2uY/9q+X46NHyA//ejyz7zz6LtW4/df3UVzGHubEx49EYijYL6ugNS+ylzXbXZEGgRVd+6DkJOX+cZ7jJbCvL6/0NaEi7WV3tj36fzLISPorui5Pcld0+jB+h8K5fAjSOATgTGGln5LpmurSM7dqqMdnvu5GnbVPGKpB1hqzRmzbp1a08ZXn3OfZT14a2UdrWV81Afx7IBsaFbXf5uulvXz/Y//CL73juVw7vvfXhj3z4l3/zf/+7f+fB/de/yDjQK34ZxzEHfLWSd9ZXjtdyZSgNs0wPfDM8MAGyb4ZXp8zpgemB6YHpgemB6YHpgemB3wcPGEVZjJ82hfwOwjWDb2KynIdkWDyCK0M5g7uK6LaBnm0d9Elr3UBz3Wa7gZ9Bu8U+i0Gi7a3DttSHHL8k16XalavVw5bR2aPxsWWmS3MJrP0i4CrwZOtfbfXcMWNFMGKnACQD27bbuwkqbV+yt4a+DU3yOgjPGVYCXqEEEQ6i1IyR7JkcVI8dnoXkGPqK/AZC4tRtoCywIdAgrXSRhVQzT3bJHDo6ephD2Ls/HhEM0TdkpqR4Cru7q/w6IaXms+ZbOZEJT2efnR+fLLvE07vX3abJwNEdvqE/T8iPDqEU/JoUN+mgSSwendisPmSd8QEAA3a+rUfWGwf9j1Jj0gbFuSYGIERtMybnDf+EljOb9GP7YQdUrepPrsPOJBJcC99GHnpELzal9LlO+yy67lK/69RsoNYnKOZ5ZFhXw/b8NozPXCM2Mw6PB+Db5lrZZI65HpwaB5tS68OqwJMeUKdrLRlVI8tKOXXGG+3oj7vRZfag6+0+Z45Jb+aYxcwt5XhxBlW2KZ6dHnPmGP7n/iw7bh98+bXluRtqvFj2Ocvvmes3AFKYJ4R7lpVL54y5PXt0b3nzd35j+cijB8sP/ft/crn98itoYF2oR9CPkm20Y0w9NvsxgD9OrHOUluET7MOnOY+Mc+9i63hPFOPzNTM4YY8ffB4uy1yOB8V7mSnogfp7rLlz3u9TQF5tc+4KNIMOU62bQeg06FP799ly2b9FCpMv/o7O8qNDQYm/CI4GW8xIq0y/WrOeCVe/c86kVI7Bdzdjo86CCG+2nOa3pfoimz/SpWCbNpzyjqgnrPzhK5Taxe72ywfQfZxtlT/FKvvZ/+Pv/p1P/cP/6++/zmp47MKAA57ytWtVV22eS8P8Oz3wTffABMi+6S6eCqYHpgemB6YHpgemB6YHpgd+Pz1AcCjcrzUAACAASURBVOZeHOK5ikbHbQRtFXzHHoK3q31tZwd9HSR6N/iTfs0jve0Wg9MOUn1uuqt1LEhQWdYZ1BJQh/5JnjTyp21o3d7bnuKrCNw2qAk0DYi3QX22fflIYF80Wz3K6u2QRsEl2wC4QDzlW2x3+5zja3s27QGzbC8giEp4EqzHHgWkKXKU5dcXOaibLDK3WBbQJX3pr3kRvIk/w6qAIbdEbe0gmA/yApjFlq1kgl2cgaSYjWLgbXpXsZYkQaANiKFcLugCXhGYgw5Q5wKMqq2OtDn+BtwAds6P65yt6/uccYVv9Ym2q6j9s0umT4EcthfNlm7LY5ulx56H8Wy9+9ft1eZ6rHXpc6/DmjvGzxooUKXAMm2zCO5Y6mno1Qc0OAcWz7mKTGhdrzzYWn3orLHaXO1mI8mba8hpm+yzaJ98YnxiTn5tUpqXX355ef6Zzy0PHjwoUFrICOBLf58xn6ePH7Jt8Xx54ZV3LHvnR2ypNNMPgZwneAAtsCVyyCK7vgeQtr884kuYO2TPXZ6TlXZ0sRx+/mz5Vz93tPyJ//A/Xp595yvL+d4B9ABDrFet79L+81nd9hXIWLYXSFUgY7IA4be/fFAusr6ex6qXT5Xn83DHar6Kx/fWkjPGzopKf5qRZ9Emn832i55hPF6t96TnbsxvdPX8RUKBoQLtzqXbai1rm8te5pw+5WbqucU3mevtGml/aZPFkZV9eQdIttu5hMYvCvt7fITPPwXZT99/685P/rW/+r98+F/+ws/xhQ7PKSPp8/zcnaPCt7yB/AeGx7NpdflxLLvGgFU2y/TAN8kDEyD7Jjl2ip0emB6YHpgemB6YHpgemB74ZnugArMrWsQMdkHHjDavJWAjQuercMZYCfQ8w9ygMABKwmDjMYOvysDYZulUwGc077lJxG45A8v+CthKf7bk2Zt40r4RyKGj9NBJ6fo1MncMJiEHiAEUGoeqa4JmCcwYNdofPQa5dJjBYZdjSnAKqGPpTKMdOqWzX74MGCkeEq8wnw2y5ZWu+m2vZzE1s2PsQ1sNCPnCCC1P2ZbwMuBk4EArnIBWBKQ7f5TTemEodw+bBRbu3r3L1rpDaJ4peQBlnTGS2L3HwhlRZjVdug1tyFQeA3VCqy1GYQMH2J+aRbZ/C0Cv9AuebPgEwk55pi8AgOG4/vHjDWzhs+gfvpeXev50vefVDDWXF7YI8GmSZ2kZyeecu/jTeSlfKyNzxt0D2eMXGwF3suaGXDOJ4nsG3/4VHMH7oRY00n27uw3MAAaivOVlTUDZmUth4k+BPK6HdllNktsFreWJP/8/e28aq+mW3fXtc8575qq6VXXrDj25527TTQgCRUEiSviSb1GEg5ACJHGCYgy2SBQEIYlEIEGQKFEUAiagyEJB+RAlQYljMHaD2kPPHnp2j7e5t8d7+051azrzec/J7/dfz37PW9VtY4jbvsPe3W89z7P32mut/d/7Ofb699r7ybgn27UNtEiUdccav/WrtJZ/pUf36ny/7gsee84b9frm8GrFuxxcx3WVkJyRGvb444+269evtRdffDFfsDyA4NqCeHzpuRf4KugpXwo9b69/5Hq7usMWy81zssh8T7EJfH6Nw/ditrqVufDjsA9d3oEkO+Jd5cuJJiedzNvx88ftEz//M+13//4/0C499gZIqM3yDaGOX3wVE332qhHxxWvfkTUoHOdx0T5hX39qwFZs6OfFEa74fkS+Z2ixrlgTzkfkpnk3+0+56ofJEM7Tu+Drhp4ix+SLdKnWiRmk0UdWpzqzJhVAr/739SA+8SOdva8tpI5D8lzC1HZL1iye2Ob8kfeVsecZvxC9mFf0aEd9M4GnrfzMOjjzzwztNGTd3Tw+Ov3o3Tu33v/f/3d/9Quf/eVfPCo6DH2xnf+VAKspXvgF0awe7fNcrePfgcD3EIH6vwLfQwND9UBgIDAQGAgMBAYCA4GBwEDge4hAjyu7CQ/p3/BHUEV8VoGiASQBY2QTLBoATr/ecflagV8FZAaaXU8FagapFRzaZ7muB5rWGTRq0r7frXQdvX+X+fWe1bWsr+uwr8Hpcl/v+0+/EvwatS7V9/uFbYP6B9q118fVbdsvhShacuzBonz3VYqnF+PlfBwBP27fvsuWsvI5+iedmStJBKcLuZR+37FUvzISEV3GQFvyayLS1BN/ex+lvZ8y1tS7GBe5K7YZki/7nnGqlxLCAR+9egi7bSHGYMbMRrLfghRCV+SQ6Vj1Z/fMmaFmcfulRRntd9l+jU3abZMItUi8SPCZ41Pnqt3fNzKIdh0+9/tuQ6vOi/X5MYv9sHjJMeUWpa9hrvqj3eoHXuB/gl+nki5crQ8Okw712GdZn+uwr1VJnXWw39zgC43qOj7M/dkJxJZnwp0dtOvbs/YQxNjDl2bt0gz8z4/ZtnfWLnNg/9Y2X7ek/xl1GxCcEsg+R5/kmgftH91tm6f77ZRzyz7zoZ9rt57+OqTZQdtwjMybdi0LLJZ8dyx9PMvtyjumxbzTx9Jl8sA/yvSfbYs1MAksPyvns2eM+dvY2MjPNTb9/UovsXMrplcJWu/NbvOnr72oz9Lr3LZ8xJcx/Qqqvrgt+YT7YzLK1NXH2q+uMO12HV2fz8r3+v6s/V7POBDnf0ooLM9OTo6+cHxy+KG/+Tf++sc/+4mP3+KTpKQInsh84+SZ+XKyf+6j9sc+5iLM1D3KQOC3EoGRQfZbifawNRAYCAwEBgIDgYHAQGAg8L1AoCLB0kyaxtkm5+uYXLLm+UchcAjU1tw6R/YPEWsCxB7wea0gkowfg22yiUIS0dOA1QyRut5PTtnHANIg0JJziaagVJ3J/sGzHGEkYYFMAlPubI9d+qpbewb33ocS4rkTP9ARJU9/NisloFdPt6sf9uvPaEGyIDGbrWTJBEnmibTIRDpN4+5nLClXftWYJHtSqK8y9QOXsmktQpMvF3g4NqYB8sFB59B1ZPQdeHHPrxdutFt37zFuxruwQ9BNvxA3qs5ZYMxVb7dOYfVSarxRyANXsSfjJWdWIQPd0I4nwiBZVWjuJTqVx173n5u6tw8EgASceERWDBR3fRzxFVEfWEvryf6xGzijXAwKb7BkbLNkKBWZ0PFVLnM/XfXJuXdrpOTOad9eR+YbSCqlSPXRD0rGzsLSH7Pfus0iNKifvtBKQ8mio8ZM3yV96Yc+159kVWCc9EeXWJgpBO4ZH/+61kAn2ZT2d77M1pNgKz+cf4kV/eCiRddtJRPVe4G82LgOJIM2NzchvMj8urfH+4JNtlbOjg/ao9e22puubbS3v+6hdn0XeQ6+b8ccVL/BAf6cTXd+yi49+rezWdu7sxeCJttnmb/trY12eAjhRubX4dGdzMf+8X778i9/pL35X/g97crr3kQK2m5b2yCbDJN1HlvST3Wa/D7Ghi/i4Blnfctvxoz8NBzGVn8vPFPOuaIpeNasMbeeXYc/hY1Yikf9XVG//cUo64LlmLPpsDnjJ+kk3oqQBRs9vY94py+Ukn/X5qyFkGluUfXvgXOu384RduS0Tsk6A3qeudJe5KJzx5qOHfvU3z37xBb1lm5XR507t2qW745Y3W6XhL6duSjP11ZdNysrJ/j2BbR+6B+97yc//bPv/6k7+YTsud5Spg9Tuop+I6WQ+o1IDpmBwD8fAoMg++fDbfQaCAwEBgIDgYHAQGAgMBB4eSLAUegrWwRzHOPdmSDCNRIaEuBRaVBn0GhJsC8ZkiA1VYs2g80u47XLeFWXpV+7vlTyjzJd3tA399isa0n1Pv1qrfeSEerN/QN+dZ1dNoHwJOt91ZeePCTs1i5BPhXqrFD8QuZBO8Fpye7ys7L9uXy8wFLferu2u68h/wy+pwDcekmV27eIlUkggTspn2gPQcl4iL8houJw9JxzIHnkyHjJmB0HPxrRwVzYwSCbrKFzDmo/J1PmDBLCjwFIBYTk0ZbyUXSBgzpSZEmm+8pOmzCa6hxvkaCo814/gVzioUgH5FGFlcJZ/ygdr67bumXMzQjrW0uVtQQjlGZOS03q+z/VXmuk13mN3olxVMb+/hyCNjJ+/PLai1vwQsZaT2VkmRG3Sbr9N3DxT0gdB6w8P+dVvlnC9QzcLZmTaMlj5Kqu2px3n/2ZEHfMFxs9e2yHg/Yv78BpHx3wNcq9ZI9dJ2PsnW+43t715htsr5xxNBxzD1Z+hfKcbcprjMezyNxqaBbV7pXLfPjhIAf1Z5xztlmSQXbml00zJ/gEqfPiN77Stra2INk22/qVh1u7dAU6hy9DMnmOyRm0BPvcle9wOVm3VmX8zJXvlWd5xZ7tqav+Iea57ePv/Rak1VI/ZfpWyws56iTKJrxPyI7UTs/2WrZpf2ixha3YdFFSuryEFrwY70Untlyb/pEsOfss6/Re/lhiLvp5cHzi4jxaX2vL+yLVkLNghY+LgiM6vk7n91/a3nn/3/qx/+lr7eiegNB8xmcaXAx6WGveu1EGAr/dCAyC7Ld7Bob9gcBAYCAwEBgIDAQGAgOB/78IVERaWuAwVraIdbcIUD0gOsEdQRutUyg4BYIGd9b3q919NjCsUm0JFBd1FzKls4Jl75OBw1WSpPRMhJUMA4VwMfVSVZ6/1O2GVDEYnVLNUBEfLvyYvKFevYaTyUKhY3wgI+WcvmWFUd4XlGuLH33KJ8eWwJVrYRNc1D0RRzRE1gBfHyRQYofnss+4VMgYhKXa0mvpvupjM+e3YUVyhWLGkGdWPccZU0boBtcqXGVLmVlm2gxRFHnmiAGveE7YVMzkqbHWOIpcEhV+mlAnX71cwQ7a8pwD+NVHVlecVraATj8zrqJTX8B1ZZ3RazJzN4VMyPuhgjWu65z7dHbCNr9LO2xTU9WEEZjki5pxRNP65TpTpuZcEmZ5bgs/ZdShnH3ECxtLJMeMbYg5s84h4W3IDu1hQ2wlUr5bKVtlM/cTfmJSBcJE34IJfqSdNucWI2Zh5uw0bAjJGqSZPSWGJLncWokH+FFb96BUprUt1M6l2UX6WBhMRiG1TskivMVW29uZrytkfJ2toeP4Xnvs4Z32B37/72mvu77DeWT0hexKxphjNRMSWyuQpX5gQtLS7cwhkOBJN7bWIdn4muUBW/748mW+8sq8bkl484XFtePb7anPfarNNrbbI297N1lprW1dvuroHXLw1O+sXa4syrgsFj6Kh23OV95ZKyliQhUFPJEp4tPawmGNtRSSMmuS+klPrvbKWnHei4iStFzOStU7qE7aiyQrbydMUeeycW2d8fegDuCvDDD1qvoEDByXc2ldsipt8J3D51NwdR2EGJ3GFKwZlFl0br3lv+B83FZZ/06oa+WUOVDXMUQl+ldPjg949dgmurFxm36funb9+s/945/+qU+e3LlzUAiduf8SdWIj6r3k5e0PS9cLGXuMMhD4XiIwCLLvJbpD90BgIDAQGAgMBAYCA4GBwPcagYpOL6yYLrPBeU2bBLAGYgZtBrRcumgRPRWgVYDZ7yMzyXnx+aLfhZFOSvR+tnif56n/4vmiW3T1zIsKUssnZf0QwIN13X4Pmo0plbWXdbG3pN/b76y7CDzVJ+ni9UG5B581Yl23yVOee1/D9RBPky5lbes+PDgWibCZmWCTzN7+IQBDtpgZQzbPmeQUY4p+lSjHs3ZlHpb9S3Cvbwb4HnYvO2B/SR+IkzlZZLPtXbXQhl9iZZaTKTEOSAKj61SP1A+EFIxEZOI7pIA+yJFp22weXTo/Jict52PN26Wd3agrMwiCCRLTPOp+zWm1+y9FIhRF/bB1z2RzzP1rpn1e9aFTA37ZsLKbuPKfjkXHsvcJdmDR6+vZ8aupMHQMlkUbbkN18cw5YLTNzRyjfe6HC6iAeot8yEWeJeYsQh+iTj8zD6XTtuAl5mI/GXT+e/2cOXc75eHd/Xa8v9eO9m6D69221Q7bm976SPsX3/O29oYb221jDULLrab4vypB5bl+WIVJg/5mbk7Q77qEnPELlhuQbPfQu8Ya2OYI/7nzJJGHjNstzQrdYgwHB7fak5/9REiyhyHKTtjquXHp0sSFFU4XvhfePjvDXPAHTFhr3mMg4xLfPtaF7ISF9Z3spCpFGYvLQc0S0b1Ez/Ts3KYgtyLJx7WKOi/mOsQlOt3a3Mm5+BHWTgIfeTr2uSr79neNFqmm3dr76Dgl4ujH2utzZ58V3uFTyOE+1mkbKMszZQ1/5e/vofMzly9tfeCpJ7706b/5Y39tz+FAELqYlPVSw+BfdRUcjvWifiEwbgYCv0UITH/tfousDTMDgYHAQGAgMBAYCAwEBgIDgd98BC4iS+PNHKeTPXeecGP8agRaQahBO48GZD3AU8Z7A8cK3IrYyBlMS772NquWCYkecIYsIDhdhViIvmQfXSgI0YKntp2bhQMRoS8ckVR1Zqokw8naKto0cDTzpAfQyfJgi5lbpSxrBKwZg4ExusNuUF99JWsmRoO6+RlnOEFKeX6R2SiRQY/9urs8BYvUiUtSqcoH7emdY07YPiGvno6JMt7XFxjBVtkpyC97nA12fMoXLEkowRecIFsL8kMCCuUdz4yDvlWwJnsTn62pefVLjBIVDID/Mrdks5glZAbZGn6vgo0atCupsQLZwh01kjcTLuoQZG1JsnmmlX51n0sDIvignD8IGbf4bZHVdXpUB9xr2t9M8gRMJbTmntNE/1pLPEsSZUGqprbMxX2kMnd41tfhPMSGctjTY+digceEE52dh+Cn31PpfZIVKIFDvaN2zOJkuZBRN+spmUCegcea4ZeMSAWzziQH8VEtjNvMsRA+5ZpSFDOQFrChk+2trDOzmeI32Eio7u/vt0N+Z54zhu69Wy+0Wy98q13n5MD3vPct7R1veqRd2Z3l7DBt8dHK9HO9e06WfpvFtQbOnqElY3dORtO5GWXgs5GD+1fb3j1IMu6PceqYc8tWjjiknu2WW2zn3GVr5ks3n2lf+MRH2/fzfAPiaWN7A9LNcbJmxBxMJNeKhPU9M4uKQWA343HdUMREn1wuvqdC4rMEbERoOGOus36dbNB1BlY4p95xqMv3w3PaojetUaKi/Jx7ybGsH8w6h3NIqvWsb8aPHP97AC6XL3rlT396kRxUv1lfjiMzbT9+sZ9758q+07riVgKstOjjajs55N0CCzPZLFkLHGLG2oKzXFlbX/dsudmzSH94fnj8kT/3Z370uS//6iccsOKq4ubCLyuDF+q89lLaIzxV1bp9sG+XH9eBwG8GAoMg+81AcegYCAwEBgIDgYHAQGAgMBB4uSAAz7JGPEkkRzHwOyXoMrj33gCxWgizuO8yCRwnuRABBpGQGRW49lAt4vmnB3IV2FVQqrx9rUv9tLXQDqknLvSabYSTra5HmX7vdeEr8vbp7db7s1jvr9tFQer9J/anfsv9JeDwrnRO4t2uYaulnxXmvW39B5rpt9C9ZE/ZYItN/es+ddu2m/VV2VJrHJp+3A4gK1LECfIjwbzbvNARMspIhYPYzQiLj44Hm53g8V4CZcUzqSY/DcJF6xyS7AySTMIDh3BumhMNak/SMOQcV/Wom18yzcQB+fKjg4JPrh2a+NZDyJh1dF/iLCtJR+gaWrRx8SU/KqKj4+pzSuYAXdqkdN/7c7dbbmFX15STfasu6esqcNtbXw/BiLroCQnn+laqyB2JOrOCeik7kiu1brtdx6Edn0PMQOZK+4RQ1HfV+u4g4zxrVyvd3zTwbJtrIiRZWJSVdsTWx709vl56wDljEC97B3fbwe1n2+XZSXvr6x9vb378art6aY3tkJBFc7byYazGBfEFwRMfJhCk8Yr04b3mDLJ1iK4T1tTmJlssWQeXV3bbfGuz3cUXx3J8dJrzyY4442xrrUiyuzefa//ks59um9uX2/r2Vpvt7ABZhcjaZXTgy0DBqGPnmOSQJp4z/ikrYaid/oMvwnIV61K4RI41mS2uyEhqWfr70/FTpz/7erXk/Z8W1CpEVNWXnP26XNfV+9u330v+xR+nWb8ytmpXrhd1SOo53dzw4zB/5kw9/mw+ZY5DfPFSMvLyb3X18PT45PO7ly995D//z/7s5z7/2U8esoRmELCqokNpVOtyUecoA4HfbgQGQfbbPQPD/kBgIDAQGAgMBAYCA4GBwD8zAstBYwVvU9BFAO9XDHvgbkhWwVxl8Rhguv+n16mnkzmdaEjQiEfdxoPPBorWGeguB3U9o0KSxaK+ClT1AUemQNi2IiVKLuTQsjyBZvzHhrRL/Ag5UsG3/S3aXrZPuhSeTYSChNNEjiC0GIv9DJAzVuJR+/esE8/OyrgIgi1mtFhODOLxxTF4laByXH0rll8wVJ9juvAJnHmmIuOOnehkTGxn2z/aa/tmkGnCH76bldL5G6vcVrgCQXYG2SWpteK2Osc1+VWyEykgx+Bk45++6JOHt6+s4QMl/oFh/HAszpGYsl4Ss+snP9vjM7o6IbXGFxOtP4PUO4Osy1cy8eESZ109fH2XM5kgfKh3zizK+puZ+mQh2y/9wU1MvXegGaO+8J+aj8K1CBllS5dDyxwxplTyHH36qK6JmOh1s5l9wTlZPtwj4vZV7rDjofLL82TvbgdfeJDIjE106FdlUyGE/blfkXRdKSfc1JnRqExciRjPk29e56yng30+nOA9Wx7379zh92JbPT7iHLH99tiVWXv9w29qj1+91K5sw6TwmQ1xDgHlmsMH/S5AfCcqI00/rbN9Y4u1wRjXNznHDDuKzzc4F+uAjLH5ZdYBpBkEmcWD/I/5+uUVtuAekcX2/FNPtCe2dtt7d3fblcf4OiYn/9c7UfOJEWcoGAYf1mLxj2JfRSKxZ2vJA4XEDSD17uAldZLjtpnBKV6VOSZwzl1wn96thV7xR1+11329g0yAfxxwYdWvedJfOUvJ+vep3ldJ1NjmmqIP3Lg6088HC6xf9eWWvlmTVJ9wyN45ZwByIhr1IMG6OjEzssbMzdkq8ohnvR+tnpx97tGHH/7Yf/NX/tIX/vE//H8PXIC2198TaMEL2GL21/rnO8VqfL+W/KgfCPxmIDAIst8MFIeOgcBAYCAwEBgIDAQGAgOB31IEDOTuLxMZQbC3vb29enx8uErwTgxXgWkC/SmAJApcBJHfqceYuyLGCgB/bVn7VkBZgaXRau+rb72t1+tytd/v+7Id+/XgVKn4Jwkx+WS7pQev9VR6I5tA3H5Fytje498QClaQ5RQbU4v3D/qwIHIQ15btylm8aqv71zO6Uucgo3cJQ2sm/0NqsS3sHmdPnSSLi3DENvrFD8iH2IFEmBmIQ5TY7nY0iU1ZmTpLTDsUfZLQCblWeiTRog9iZnVmlpGBffmujxyS1OaxSX+ePVMp2+gmP8yokT5wy96KHw6Yxlt+kEHmVreD47ZzdZvterhwr/ATJzNsBEZyKjdxsRNZheUF0biEkbjx07/ggC/ed9wkuRxx6rjp4+ntNKX4HBmeSgbiSD08PyhrvaW8QLfjT0XpWGc8yvhmSbIAEhQJawGi10P3xcz2rseuTqlzJCGnfb8uebjPlyX5zSE6j/busbXx2+B3t12GwLp+aaO94ZGH27XddbY9rrCdkq2rjFQuWf0hTaf5UH//OIX1yeLi6rI4JVtwBpE5P+HA/nXISUjCI86h2yArDDXx8fLVh9ra3XtkPR23Uwi70/17kGTb7e6tvfbNJz7Xbrzh9W2DDLJdzsNzu2J/xyRKxU4iLtuGxaJjhU9F5FEHY9yx8Npxjd/TvHjfZfp8RHZq72T9cl3vo8n4QYVrcDr7C9Kx1kzXq/zyGvJ5uXTdy3XL931teT1mPTN6FPJeMi+enyhhrQ6/Jqol3mmSdKEjqWN1fAsG7QNPfPlLH/g//re/83T2jzsB5PghswzJsslxPxB42SAwCLKXzVQMRwYCA4GBwEBgIDAQGAgMBH4jCBgkJsibhAlNiRwhJLwhir1+49r6/Oxo3XjNL+tN8hyFdUbi0BJxZMSZYscLMsKqhY1JZjn4lBDqz12u+hRJ19ussyzMcG9bfga73Ft8VubBfh6qXaV8SxYNFffbLALQul6S5eGGJ+ruD5TLtplElpBVXD1/yiKnEx8g5ArLiRRDPHq6v8hqbmGT+549U76pbYl085GS7Xp09NDvuxAlZh+pyOyeXPVDp5L5xXlPHt4/ZbVIltCy8DkOmLGlI9bbTsZWZjJ+0kZw75cDzejxxKUQbG7ZTCYc7Rz8DiL4joJJD97QrkK1ep+gvzKkyH4y60zSR/rr6pVL2W55EjtFRPnlSYk1iY7FeVnY9hwu+1i0qtf5YbeoO/GpzKdgSX3JQ37Qv9ZIkVPq8CugzgmDwvXpfVhcq66v9STJ0RbWiWudjWWfaRsxnmStMObSVR751cOsQbKH+jl5trtlMhg6V4zLzLIiy7wl24hns/c8FN8tjwd37rV9vlZ596Wb0CT7bRvS8vLlWXv0oZ12DYLs+pUtDuM/48wx9EmsoSPu8q6GluGaIvFpYf1YfH/ExS3LEkbxKW3IzdY5op/zshpZfxueXRZqL2tOggyE2p27e21+OG8PX9ptz9692b78qV9pO5evtC2eV1d3WZfOEAUG7AwSSjyTxUiV8yvRanFl6odntlnyDvV15VwzGOdKIs13QCItcxdZx1SksHKWmuuL+/5cevscaW86Uyxn2blgS29QQpc1qfVenHxHuA9RTsPimfkqYq7WsD5IvsGBRubw6CTP+hkSkvdAPXsne15BHGITemx1c3MPSD73ukcf+eDf+9//7qfovc9LPE0eJ5vBuvcxaGOUgcDLEYFBkL0cZ2X4NBAYCAwEBgIDgYHAQGAg8GsicH+QlfiLaNL/rrU3/47fOXv00Ud35ycnu2S9wDFUJkgCVKK36ltBa9djsLd83w13gsH2HkzatixrveVBHf15+bp8X8SMflRga5tF3V3O5wTlXHu7m9+8778H5S+e7UMQOf+yIQAAIABJREFULeslETWVrqeTNFb38TwoE0jFpjdwTX98tNgvfZWZ7rt+/V5kw0wkQTpFaWs3b97K+U5dj+SNW+QYMNNYgXqIIvFw3sBZn0PymDo0yeIRjpTm7kueJCvwKxldkCV9LNbpl884XR2p0++MAfJnhUPGcoB+Y2sldvMlP/SFooO8kQiZnxy3G9ceihqVSKPlOuGgDT8QYJGwtHSMlu+zxqa2vt5sXy7207/4SIMH//fSdWadIGORsOjj8blk6mp9r/PabbrvLU024++iv3aFnTmoTCkIQsbmhxdO3KLKXPgOaMNxSoyZYXTsWWO3b0GM3WkH95jrw3ttnS2Vl3Zm7TrE2OWt1XZ9Z7PtkEW2AQEH1cPA1CO+Th1zkAzDen/VL8qW7pvXuhcPOrGG/ECCWV4r/NjUB6FTxBZ/DzLvGS+0me1mmB2ZSXZwu+2ub7UXn36yfevJN7Qbb3xj22TNRBYdpkiFfOPvy7mk6jQfuYJ2+eY8dwKq1tJqiLDyOdjFezwFM3VnHdK//w1xfI6nF/VmHSH73Ypu5Z2YGtWTTD+eu0/q635lPJNO6yU/lcs7Qh8/5tFtmjnm1srj42O2oZKJqb8M5exgH3kIxtXVOX9b3FfJ1J3PVlY3j9fXVj9//cb1D331qa98+if+3v95b40sPrhi/wBlwaq75qsw+W5jGnUDgd9uBAZB9ts9A8P+QGAgMBAYCAwEBgIDgYHAPxcCU5hVESXB1x/+d3+w/ch//GfX7+wfXz44Orp8d29vtrmx3S7tbhNLrhLnT4FmDxpRYJBZwbXZKlUMBnvQ2gNW63LAPXaIcCdJbqcg0+DPn6X36c/2rfvJY8Layg6rZ7e2eSbRaqX6RH9tLSudIYjQPUNO3Qv9uOF2tyrJkSJWJWSmqmQchwQBFZriPn7w7H+kUopagDCimFFkP6QiFymeVzPmKA0u4qQez/HKCLgPPuiscUoiqHmyp051UOIXCp55/nme1FR6M8YQLhf+S8z4ZcX0RccaW7o8W2wFQmXSpkqdubgqbzxu5qBkl0RJMtKwlQwf2hRHTzKRyMRyX2C2FwpJDoKnjv8Gi7hnA1XoXoXAOTs5bOdkz7zjrW8MmSMhVWSHrtBO51W2dZ5L5KUj/Vw/9BcV/1V39IsjdSJR8lW/sE87oveV3s9K7y334Ts9a7OymrCPnDJZ1yEPEUpXrUPmTXpsd23602U/RGA/CTG/PGo7qAKfc2uyHx9DqOXD2WyQUPyO7pExBim2/9JLIcZ2Z/O2fWm1PbRzJV+mvMyXJXc5a2wT3a5ANqY6gMytK8ovk8b2NBerZodqlYwpi0tL29luqa9o0EfrAznXFTLGZhCdkq1QPfRabbv4sL92D+KSrZbUH0vk4fx8/6TtHd5px3z18qkvfqa96R3vao/v7PJ9CL5qmSwtekN2HrvdV/uMX/uZmNywlKxzqyOLdnFGXkTwIWvWMeg3WDO44EyvE9qyXNHjmX1ZJ+jo68OrSzVzwHxltUzPrjS8X+BRvGnN80WWq8/TOxT7Ol7FNZsfVZJkZuT5fHR40g4gMyWGzb50O6314qXf0zo652MIpxsbGxz75tdhz14gy/Ajd27e/NB/9KN/4tvPffsbGHGllPvdpn1HGQi8nBEYBNnLeXaGbwOBgcBAYCAwEBgIDARegwgsEwC/weEn1P9X/tV/rT386KObt578+jUyHx7iMO61k+P5mQEcAXF2NKq7DtEmcEW5v5waTX0vFYwWUWFAaNBqXa9fDvF6wPegz9YbhC+XLrN8XW73vvSVra7ba/chATRyeZZtMVyP7/iPY9abQdNL2SpCxsH6LIHT+0h89NJt+Fzt1VI6lkc96Zkw+bXke7/us89muGjxpVt3IDEIRcyyoj5jdRz8vCyKD/TpuqxfyHKf+hCAk3+QDJJjAAFxgCWznbChXBWpKH6yiMUk8sw8hZSA6kKuMr74Wp8km+csSWJkGxt9uF8nHeiILJo3v+HxdsrB70UaoGKy0H2VzPC+Pwdfnlexq7eZV3r5JEGYyqnePpISfTuhso7HDW3SgxIa1kmQLuNrnfO/HlJJG2RkZR2WL5OL6es4u3/WhyRLXeFqNpZOKXM6kSOOFS8yZs8ZCynE9Qyi7GhvH3LlHueL7XMA/0G7vtXaFgffb85O2yak8qXtWdsAO7hDMHTbI7oFAp2SSpJMFl7V+8aEQPy1rY/Ve9wK+STOy++p/vbZQBNLjIP3weAAOxt8dRSGs63zgYUrV66ohkypl9qMbYSc899e+NZX27ee+nK79vjr2trmNnanj0eoEb3accZiXDaOOr+0ObnOPYgxJ86DfscX19lUJKElrK3PPfPj+5C5RMy3wy2qWSvo8G+TW6tPsbHmuuHZn6b9O+Z9v+oENXFFPy22q9W11LFb6GANKZd3Ul3IuH34gA8XuIaO2eJsu3WSZN6fylijcJ10MfRsa5HbOyvz049c2tr4uf/kT//I5576yhf3qQcKBiJLNspA4BWEwCDIXkGTNVwdCAwEBgIDgYHAQGAg8FpBoAJI46tfpyTuJF4z84qA86WXXuQLdfucPXZ+CYJs18Buf+/wbHdnZ2WLwJhMFPggSY8KWBO8ot6nqrmwFftEoean9AwMg9dlSQPGrsOgs2QvfLbuu5WLer8LRyhpgG2BRGAYkAWSXATGVWsDPhBu02a7Rdtm+XT7da5Q2attm8hO5o3P4x/jtl8vlc2iwvsJwIwdg+mDjd4nWVYQOX3cZrRZ9LXGJJliTdXrc/dPgsIAfba+yRfwWnvx1m0Fi/ThIPwqdFjo8rb7ajYW8xa1E2lk7N2bHSdtJkadewYVdnI+FZlj52wTayscKn5WJJmiKRJS9hdkgTLzTIcXv8JklTC/++FY/NWWtLP2hsceydbAI7cVuhb4SXqgpHTljLNSaT/nT/19CiSCotMPKuBLja/mWR0s2MgrY0Zaz9QqrNHFAJIhR9+QYNO6tmUhs7TWXVHOge9Azal+arevI8iO9SJ1hUVSpc99qA4VU/wSpRgUccJ1/5Ctinc50g2SCZ8u7a60jd2ttikJdnYEGbbW1jl3bM1BMvi1GZ44X4xbQkn8QwrJnNG/CD3HwPzhoJl1vlv6aXFukxGHriKQagwOxvouN+NsuxCJGDuH4NnY3GJ8kGXYU8Y2l4EfizhirJKee3tH7YnPfqo9/n1vb2+9/ggkEdsJ18kkw3WnNvi519DpEbz6b/zSV9uz9qhPhzjMrbLOV01p7Lu2QsainNWR+6wfhELaU6ufWVv0l/yy6K/63PppW3xLE3WMwz6296v36s2HFezH/Mcf+6btnHeSNXHCtlOuvhQnkGS2ebabelZXTzlT7tgsyrOtrY1T6rfWyNCDHDtC4S/w/BN//j/9Mx///Oc+yYutp3wGg8IcDoIsszb+eaUgMAiyV8pMDT8HAgOBgcBAYCAwEBgIDAR+bQQI5gxOOVeIXWWrs9PT+eycLJrj+REttYVonQDc4NuMC8moBIcVc1fAiJw6LAkgZV2me58NFJfLsmy19fYKZEvHFLxPeuxvPwPbIgcgNwyCqbd3fIrH3CtMiSx9uj3rtNf9iW9hemwpHGK7K7Castwnz7Zra4lEsb77oHyC8z5urtGrEMW2lKk9fkwypaPGWmb8tzB3V+Ot28TRkFkhMcSCQPwMQpNBlk9Ia99eK2QAnbtNkvtVMrrO5kfW8rP1opi5Y5Eg9KB8E6AWRAP1EnwSKG7hi26v2FO36ngKUbbAQ4LmtLLK1MtBS8necrPuxuZGe/yxy+3s7m0woT9jEI/C536/MFZEDtWxC+YSXt3/XrfAdvJvGfu6t0+oq/vnhdoFVvTtZKR1rpkcmg/DtQZRdeEjnaZ+XsWF2eCuxiCrYXZYlqLviuvKOirEa84WvAO2Uh4f7beV48O2BSaXNmccwL/GuWJk2YHFOnvuVvn64cq5BCXz4bgw4XrXTsYv7jA8HnhfhOH94alj8Bf5yDpWSWvmBlIzbeKZcdZ67DhK8C0woF1i7/wE0mcD8o4+l6aswF0+JPAQ55Hd4mMC6/hy89lvJYvsre95T8j0rD2yELOW4kv9LdAry3fME0CVz4VXSU1zJH78LF4X/nGvHqRydTz+kkVIrfd97jIbkIbzbPms+q5v+aq8JGD+5oGF9krHRHzS3v2MncmmxNsOX/O0ryU+8lJ5vXx512WwNQu5e74H2fjBnfX1//u//q/+y5/7wqd+5WleIJozD/Dm46uV4jfKKwuB+/8CvbJ8H94OBAYCA4GBwEBgIDAQGAi8lhF4gIdYXyPTg5hzbW19fjI/nUOWEZOvrZA1ws40iAIC/Ry4LWZm7eRaABr8JWAlU8VgUbLFDJHUE4y6zakC2JJP18k+YiU3yZs5Yr9Fob0HxVVfAT0Rvh3ROwX4KqIYgcYuBIDBbe7Vrdyy2i4/Bc8heWK3gvCF7OTLsv/RiaH4hZ6MXQICWcmHnFuWAFqfpow25CQ3Qkboz2TXPpZ+vQjsDcj7Fr+yNeNQ9rvH83bvgHO80Gtmkhl9SHLDf7GJNzICPNacoJj/SlCIl+yDCClPvfNaxjGQAdRYwC1FUexke6IknJgxl9l+KZFm+o3+ozNnjKkPH8qmHuCDTlJcPzO+lDk/OGnf/663t4d2G19CrEPlyZdJH4k5JylYuMZij/5czbRTn8yop0fRQa35xU1r1BN7hTWepOAqLpY/IVbRpe5s12OonsclPOdeqbeoKzIQkZJ6eLCwaJsZXAUeJiUJHbt9NYAPEmo+C8ccsmTONktJk729uyHHzk8lxubtyi7nia3O2aJ42rbxcUbm2Bq/Fb4WGad0hnqzJVVfSUWu7VpLzmEKA/DsLN817aIp12xhVMDdfQLBfyVi1tDJG80z8hOc6Ud7xo4PlnPGmfHKmK6jd2UjXx+VDNsxOw0szCy7x4H9z996ph3uz9uXPvWp9jt/z7/cLr/uTe3I+cAfs6nyDmWKPDut/M5h9DhVZ425XnSR5z6p+GC/em94MMuREqwdr2uetZssLzIefQN8bxxjiDHsmP1lrzkYnEZee64fyEoM2sc5i05wSaFdncfoLDyLxJWQTJYbeOR/LEB4trFZOED8+rdRfz2g3yvnjKnOt4sENf6HBwhP/LrJmWnvv37lyv/zP/+Nv/bhL3z645Bj6IV+xntFBT8zZedRBgKvFAQGQfZKmanh50BgIDAQGAgMBAYCA4HXEAIJ9H7j400g9tijr3Mb2pqB7NWrV+dr65vrMw7aDsk06TLg8/lB/QbJlgSS3EvPGOT20uUTeBvlUxK8oq/3tc77ZRnrDFLr0OzKaNFSt2P7g/LWdXs9sNaWchUwT4Hwwmf12qsCb/tEJwHzg7r7s/q7Dess/bnfW2ubHxDoZVmmy4V8+i46ui3lvJcg8aN3+3sH7YCvHEqalD7GhomFlWmsElM5pyzsR3mgvGTZOcQMneljHM64MyfTuKlJxpJEj1lEZDLxnT3ukZ3IgxW232mPvBiukFpTtlG2u0rYIC7ZlW2l6Bd3iZ0iF+bt+zh/zCQwSRHxzrpShnFeED4XPtedbmK11Idx8Fmb9CobGUfhVfMyzZN+T30lcLXnurJ0nCWWJDAL08mWA5lKl1tcxSckmThKaUxreVo3+mSdpNic7YenZFrt37vdDu+5nfK0Xd0kW2ydbCO2T66TjbXJJEIv85MhAiu0ms3nhxUsWnG+3OLnO+gPlyn66DyW752gtAWAFwSlJJ8EUbhPcUeb5Rxyrm64ByM/TOC1E5sSVRLj2VrN1WxFz3Jbn+Z87tbQ0+127drltvPt59oLd++1bzz5pfbUl361vefqtbbKxwUkpTy0XoyL6Kw5EEvbLGYYFvYXmFtvnXL9l/5Lz8pkPoUN2Xxog2vVi0ytL4aBD5BdmWNseM94QkeJ3zRvfX2EALXP5J9zop38LWHu+5oTC+3m7yS6XRPO+azmyF2VZo/B2c3XKnNv7UWW+s9vrK7+X3/1L/+l9//iB3/hJjm6WmKG4nc57wBGGQi8whAYBNkrbMKGuwOBgcBAYCAwEBgIDAReCwgYTFaw+euN1pBRnsFQuTKt1vmm2un5fHblysqqX7C0dEIsWRiJyCtgdcuXNswMQg0BYxEhBpGWkCK064tl2adeZ32XI3MtwX9kCUBzdlL6Gi9WzJgxTfYMZPXNEmJlCor7uCuzyrapf8gGyAWyXRJQL3ybCAFjW+qSLacuCagov993q5bHQnKKNRAL+AxZE0wmXwyivVVefyM54dGfzUzK1yUlWygL/yc5dfesFMnLW7duQZBxnhGR/QyWqfJNdAI5s53EX6PoMzPK+zlZZ1IF8VvCRcII/cEmXSVAtI8Ml8UYvIeQWTmDEAsRhU4zgSAA7F8AIcS6MIMs2T3Wqxu7ZhG6urynNl91RLK9861vwSe37hZe+uXPNSCJYFEeT3O1Td9SGNcqTjo7saEtfuLQ7dozWxLTu+qjjNu5Y4oirvgVnNBHddaiWWWxi06XTn7iRYmfrs2p3nVUBF21zdTNG+XcniLk+Pw65fHBXju4Aw8yP2xX1sm8khiDmNrgfDeJsRlreoMf+XXBUQzMUrL0TDRtu4Q2NytbKe8l8kUySvbU/ELDxE/P6LJPxoO+YCVqzlPKxbvpo+Ps73SaHT8/x1i2q1/WCbdutbRs8MXKbWw//rpH2x2yyL717Ofbc8890z78/n/Ubrzuje3Rd77XPyIhjdSTH2vtbHqP6Zo68bKtT1m92cw69h3rmWeXUczy63pSwT9pBwtpJuUZLbhoq9aSpOEpz0LK37feLXNVW2insWG+CEnXwGSPTv6NOnPdQRSHIOvj4LqaL3UWRrZJSs5y7pr2yL/LxJzNVjmfbmO2+s35yekHOc3x70OOfeQXP/izN0kVZFBZvXQ29a18WTiZlenTg/UXEuNuIPByQWAQZC+XmRh+DAQGAgOBgcBAYCAwEBgILBBI4L94+nVvKgpEhD4zsjguE1jvEnDy+cFsBaqglXbJGYM0s7kSaVafCqoJLA0+E0xTb/mn+WC7gW6Xs2+vs3+C5enaZazv951YS0YIffEqbQlSl+67DcNLD8aPj1wRpqZKZLiNTgih71a6XduW77Wr7l6nLn/a6cU26yzLct4bYJtBojvLcvbvY7SnU7LGGWI3+YKlqiUFJAKS6WPnSX8fX5EdEDiyKvqkOyiqsUI/OM50Yw4khdzeyBcTo3zFg+i9Z3uYA5yCc7kFA30coxqisVTSF0UBwis/SRh8cm5k3FbZludYioSZt8cfuQ5xpN6IpS1+0if+Tdect6Vvjg8SN8QROgundM8/1V74xc4kY6MZPr3or8WvGirnz5K5iY085rm3WeO9uGpHDHwF+rNZUVCsBROywR93jzlb7IRMv3u3b3E+3H5bOztslzZW2y4s2gaH7/tlynVIsnWuboP0EH5JsXzxU6NAV+Ny9mtN+RGA5XUkOSfcZhYWJshOY1JF77+MadXVmK2vc+ZiIfL965yujXA74JfzusweQ7f9vXIiWdbN2vqsbW5vZ9yPPnqj3bj+UHv2pW+2r3/ly+2pL3+hPfKWd+Cz23P1bRaSSd/612JDdU7Ydz/TnsXKetC++NJ9eeze+9MXCUmv/rJ1ki2vsQepJZ4Zs4Tx0rro84dTWOJdIhMuRUyW373p2b6e+SehXX8LC1/fwxB09Ik/PHNlsdTawv7M92Nztvns+mz1wzRwIP+f+4WPf/TDz/re45yryQXel2f5Mf4dCLwCERgE2Stw0obLA4GBwEBgIDAQGAgMBF7NCBgMLgeC3znWBG5G3QZlhqZe/craZc4cuwZBdpkAkVidYJ0UJIN29eXMomRlGFTDElBmBPux5wPB6X2BJVUJTKcAUxGfDWK9ph9tFvWXG0V+8MVMnIpbpYPW3k95i0kXBqsJTiUKZC3QU4OSsCCA9sHYc7KTCJRA1j4do351C5qdDay7b+XXlH0z+a3tjBP9BLt6EmKj2+hb9wy8GSaZZUhkvDXWnumDy/REgOAeT9GhXeoQM+CfYQ9DPKOHcUpYyVE+/+1n29wD+SEOPHA9/pN4sspB6N7LVYU047yv6BWTafz6XvII1YMe6GDmbxVccp4WhEFIrjWdxEuDf8cPG5OZL7YCmWhZ/BMZhxngp2rIsp5luMkZaqsb6+3RR67xQQgzrMhOm/SLUVg8fY2/hRcUCM/dUH3NU83OQchaZqHWht1q7mwXm1zFtT9rC3/C4XGvfF9XWlNnCI9prlfI0FtlApNVZJIP45J4NJsp2/NYW2tiJNLUu4VU2ZPDg7bHhxSOD+62s+P9fJHyyjaH8JPdtQ4R4wH8mzhh1qFeZqQOX9xCSNV4zYL0HTOvCPWR9O1Nlp2iVJ67wNBi5qP+14RShR/KnaDD8drftRVjaVOPMtM7SUfHIBOFOGL+yxTz2dT45XrGEeXN9lr0E2dIwq1Ll9uN+Vp785sea1/95tPt5ksvtM998hPtPb/397VLj220UzFjLHO+MhE72sCer626LL4bFudE4s71a5tykridzLOu/5Tv7V5n+DJnvUj0nZCmePE+sg6p66WwKFDmvFvOe/zQJ359LSzbCb74dMoXK9l/Hsy7Ps/Xix+sE/4WYersDFegD9fabGvz9ubaxscuba3/wz/5Qz/6sY9/9OefzTtS5JgvOkzZVJwjy8LVwqQqx78DgZc3Av59GmUgMBAYCAwEBgIDgYHAQGAg8LJCIIHeb8wjoy9+qzMC++tcHiX4v2KAalaKxaAvgV8PVAm6l+uU6fY68dTbvVqWr8r6rA2vPlfgeb+tdJz6KvegTNfRbXe9mlT3cnmwf++zLGNdr+9+dZ0PyvV2SQhLf/ZqWe4nsRXd0mnT2LuMV/v0/r2+B+vKL3CCINje4WB7vhbojNGzSKt8ja/GHPuLwHryywwy9PSiTgzyKwIpmiAHlEkWF3otEkEldzFGCTTlVoj8Mx/cS+CVXI2bhvgXsgzbHGrHlxtP0Go2G1sKIRIukXEkiaS/fa76lOmfBOHyfJtltyy7jIu+dhIkY7OCEizqdhpRYeRZWBJzXbZfzQrSl9CK05yow/aFL5AdPvefB+WnkDC0JmGH33sv3Wy3X/h2O7z9fFs5vN0uz+bt2hZfMOTKqNlKyXljHIA/g8Rhq10IVClQKKGo0tbyexTbJiRhVwJR0qsIMt/DiTzKVNU6moY8Xeo9kNtTjwRTxoO9PoYun3rHEBnsQCS6drWRvvbnp5zzo480ckD/ZlvfZDs2iVB+vfH1jz/Wrl/mCwynR+0rX/xCe/rJJ9oa88/yxb64F6Yh4tBlNp8ZYtHbr+jvxa+mWi5WcM2t8pb+fniNT9b5btCv/C1Sr/tuvwd/9l2WVY/roa852322vv+03ddHt0XVOR8sgI9mXUOO6QfPd3c21j92eXvjp370h3/oAx/70M99w3cBtg5x/4BckGP2G2Ug8EpGYGSQvZJnb/g+EBgIDAQGAgOBgcBA4DWJQAJxIrEEzwRouW6cnJw8TPj7GFkzl89PzIyZSJApZqssIACzBwGjQWYPEH3uQaLXyuwh+8RskSnNyOBcOUsPbpXtunrQ2nUty3jf+64SiPtslojBvIGtWrMVi8Daa48zlStfHK5hKRk8E7nTQ/BzSBvHej6fBgoJoV9o1NWFr90fM820Wc2Or/crvwSo7Ne1huwZSHiJqElCKZArZrlgII/JaOGuEDJ0vrBvdpB6+KAeX7DcRwlWrbCvOnjWJ8dRvne/1Y/SyYaGcli+h+5jvxJ2pGfUoeUiwNSX8dJP3BPKT76veu6ZOCujD55Hpn6eOxRlhzoxJ/7vmYYSBlvk1OzytT8PrddGzZFjNaOKDCOcylzrN8VZq6symrmwU3NSvlY23dQeyYv7kkMh9hb4oEfNjDhF0sk2bV/4RBP4Ouea9euIHtquJw59nay9rD/qjw8O2t0Xn+MLlXfaClsqL0GCbbFDdXeLr1SSZbaGDNL5SqX6JNRYSQ4QE6fJ8ipPdLP8DMb9Xv9gulw//V1QrsaGX+FB6Ue6mHVmYdq/sr+wxX0d4F+4OIfZwqrRjKlwdilkPTBuMwYvsrYKG3fP1vzgD13LhiiCG2TtY9eute9/x1vbV771QrsNHp/+pY+117/57W37dW8JsaZfwT0vYM0J1Bs2XR3OCcCGOKx5tRaplLzL+kWFX7/s4+/z5vqX2Pf8tTMIOrMwTwSGv0HKWPLucnVbZQqyNuXMQvTmy6bOt1hPfbTjfeba1wSPPJOs//2xTeKPDwhQjs7wg4QyttLOZnfIaPswX6v8iT/2b//Az/3Kxz78VUfDf5x1NLEoFsXxlO5FVW5ikLtpfu5vHE8DgZcVAn21vqycGs4MBAYCA4GBwEBgIDAQGAgMBP4pCBgtLv3/squb12488hgkmb9tg8ciDMLS8Am2KTgjOO1Bo/oNHPu139dzZW0YrCvfA/oum07TP/bzp5y/nj3U9XXb3e6D8uruJFg/byoyBr3oe7DYtuyPW9q0YYj+3eR7f/vZ3j8e4H2ypAikDe4t6uk6lm2YIVPZPxB7jpe+Xdarur324rPFbWW5ahs/+b4AB6A/R1VlMiXjyzHy327PbWqVZVS4RoF+q5Pp9AuUZvv0ehxmHP7v/tRpR+ZH8kCZ3k9h2uJnMTGOiC4xTOIh/dVvFQRkilhYNY1LomN+chxyjF2W4FhZXOKl7+r21/FTR3yOsvqnP/drb7LPcp33HU/buk4JwcL7os427bvuutzy1bblZ22GiGE8ybZiTCf799qtZ7/Zju681NZPD9oOWWJmjV31zDEP4z8nc4zzpmYcyr/CFss1yC7ZSbdksiIWvmtHAterv2Xb2pVsdB1VKbynh9QvyDGaag2ou7LxxESdXs0OW5BjKEgd9ZVZh2/JSsQ3zvLqRdwK01pfhWP50P31urm53t58+YgxAAAgAElEQVT0xte361d2If1O21NkkT379a+1Fc5kc7zRwdpyWfiF12hgXXYiLvlk+HKyzB1NTuinRTvly4XvYmXpmLnV0nu3sbok+xitq980j9OzJG5liYm9/wMBfwUh3Hrm2AZkqD/79uKa8RndyRxbm/HtS14AupIpuXa4tTn7+O7m+k/+sT/6h98HOfYVNmcyXuevcvocxygDgVcTAiOD7NU0m2MsA4GBwEBgIDAQGAgMBF5bCFR0li1ya5sEgo8QdD7KQf2bx9OuH55JqDDoIyiVNOFa264I3itWDWIGejlbiycPpM72vCnj4WTKzOGA6gSpZmoY3GZb3FLAuxz89vvIIa+jHNtU/XtQGZ6AFnToSjJbjEwp+mPgan9ZGr/WWLxC3Vvfg1NGF3JMrke6osbitfzt+sxQCukQExUkG+auQlzpb+lUxrHxTPacw0vmDkqM9+MHhsyS6vU4qsNku0wkD3aTocVYCsca9/qGB523dvMmX0N0XL2YNYaOnJOFXqRlCdIaHOOEdfjGCGt8TiXPOtWzzjKHjqUU23eVJJczgWXqgVBKaMJ0Mo5MSEIJFbdsSsZkNgCG/8Y+2Yin2nHcyO1usyWPNrFz6ZllKNEQWeeNjrpQGT3ObRFUZlmpc87VMSwygCZXKlOqMEw7Mn2efXY9iJEEp/CZZRSiK+QJ2VS0SxBtcBB+Mt4cCWtDnlBM4iNklnKuFMmxU7LGDu7c4fdiWzvaazvnx9QftytkjW2Tpec2yo0sLLPiao04zxZ9yoAYoX5oCM+Cgwl+eT8mQjqyZpnJ9Fj0iXFYP01X3kfXZ5yl3rasf0GbihhnHm3Hlu3a6e9KXV23zJV9mKBV5j/98Nt3Xxvl+xQKO/eSpujzK498CLfd4LD+d7/rbe3eZ77EmXnPtC999rPtde/4/rZ6+RpSM+ZBoqgwoHfG4+hDOOEbBmKTT0Xw3tea6MPIfLgqvLHS95tx+cVUsQ1JzjvJLLYDvt56DraOc3olVJ21Z6ZYztyjLTgyzhmyzkXGFyjVDdm1scmZeUepTxt9/eCHeB27fZTJ1QPW4BpZY2QWruxtzWaf5DS0f/iD/84f+flP/crHvjb5qXUmsf7AZs07/pSld7pX/br19wmNh4HAywKBQZC9LKZhODEQGAgMBAYCA4GBwEBgIPDPiACBGtGlpAbR9rt+1+/euPHoI48QsN0gg2zDQNVAkJ8BHUFipyO4pyoBqU0U7yVelot1du3Xfm9AGZW9H3KeCWVd/6nHfr10HcvXLtN19av8kFk0y+2Tm11dguVuS52MqOJs4Fi2EbKBXtZVkeCQWClfTx0yTV4kiSRM1Kt4JyHSz7HlhhB6itKLuDHAn/Cjk1a01bH3ftmfNbK85KpuvQhBhlXS+jIXGnTrXIJ97onyaYZ0gaw4O8WfAFA+R2cnBGTbGIsFbRjn57P+ui64nvllv3MIgxBcEnSsC8aQzDacMXPs7PQYGVGghCTjPmqQ02FZMPp7VtXx4WG7vHPNpL3gZZc+xnRSBXatK3Kn2pUrzFCMck8Km6Oz46l83dccXTyXvq5TPf1emfpVXZYBEyfRZr3jXC7WZaur9hnvyf4+54291E73brOl8oDD9484X+ykcdZUtlb6dco11qJbeCW8GEnWjnf6kHUqSyj7mFXEvzy6zVSiEaHIuehco5Kl8WtxLf/6eDpxXaawqyFKcKtbVU5jdoyhwGhxnosk8nqB6TSnSMQuj/XlyZob3wPls2WXcXLWVvruQSTt7u62t33f69sXvvgVtkKftaee+GL7fbdfajucVXbOFltYtIzHrDGXodsZHaXFbZ3lA7PMmlyR9Eam+6YvKdNYHJOkltlu9uPzIsn6Us5sPAs0/2LcISNZgJFFprZk8v7ilnUdT6ffv3rqcWvtxsZGMIPPlZ+sucGxZKplgs/4oOca2ypXD/igySfv3rn5k//hv//v/fSTX/78E2Hn4/eD2yrj3vhnIPCqQWAQZK+aqRwDGQgMBAYCA4GBwEBgIPCaQoC4MqFk+6P/wZ9of+bP/4WN46Oz6/uHp9ePj4/XJTXMHIMkSCoJYapRbIJCM7mSDWFkSyF8pJV2itTFSlK16Jagm4wMw3sJGyNOioRNAloCRrOt+vlUCcL1ClljyX4Gl0RQCJi0SRVUMZjtwXLuF+cMFZEwiV1c6L9cet9ut7cZiPeSIPrBZ8Z3TjbPWshFJSc/0K8uCY6zYFBarPM/EiKLIB+ZPo5uKyMTZogw5SSRUiStGOuMLBY4GX78I0bxC8TZr6iuZb/tnK98CqT9w4WI4wWJx0RVkA8JESyUS+jfDfNk9k3YPr1je+AaJMGEY7bzTSSVBETja4f6qd4UTJvNo5+6YfaY53A9+vBVDrO3Dn+46ncwUl4MOzL4k2ewzPa7KWOoiCLwyapjQx6MRUgPjKqnZ1nZ159jyPgmItYtje6Bq6PhzVyb2vFnc3MzusiizBAkK/EKnaxZxrbOePyC6MHdO+3wpefb+cG9drZ3h0P35xB/M4ixWbvE0eyrZI7B2OTQfgwEF1HRH1gfPeWHDc4pq7H75pT/aXWe+DlkCbtQaJA92WJJ33rfai7zPlIj9tHlfFEybV5pmqqYi9LLauG/euRdcrhKHuE5hJ56qjWSJcc86eMp8+icFXHFmlaQNZQ/FeA1g/wyE+8Nr3+8veMtb2xfe+alduuFb7VvPvnl9q5rD7vRlHG5nXGDPhKdPSOwxmrWHuozbp2PL8iJR309d1oXPFsyJuRAPc/ywyGM6SNp51FfmUfmMO+zeCivTq7RIdb8sq0StG1z5MGTswlXJIIlkJGf4Zx/s/gfEsSBoSTrbNWvWELIHUGYffZo7+7P/Ok/9cPv+9qTX/ycSwnVGnIaXVDlODejDARebQgMguzVNqNjPAOBgcBAYCAwEBgIDAReOwgkOvw3/uAPtCtXr29961vPXIf8uEbQSAzo3soEnMSlUyA6hXUSYhXi9eB1OcgkiOYxWwkJJg1AJby8dj11XpjxvPqnoD66DYwhPiA0DGhXJZEWtiuAzTO6LL1toVu7yKu3t0WQ2NS6IhXKru1d1tA1ZAKO936ls85uqq2VPaZl7IzfdjHwmoP2y9A0zqk9IJWchIvbxazqdrstyZ/SU/0M7st+ZfMUNATtEAp3D47b/r09BsHnLMFVsMXMbKc+7k5gdTvheJBxTlCsA5O3uuPgfWQunDjLcrv3E97WS9ZoC21T1k80lAz1i/5TH31Q3kyyuQQa2WaPPvIwWWeQMNQ5zuWxZyy6ZD2mzyCtFhldECe1ZsqMMhkB18Kg/K/MqCI/tF86J3KEHj67vsyC6/bV6HorndhnKNWG/46Z8XLePudoHXMQ//Pt4NaLbfWIr4ke3mtXPGdsa9a24WK22DvKprsQY6uScA6CvmK/BpEix+KzZeKnkC8/nE9tusLSbZqPM52ZitlONa9OU+mxyftscRY336loqTGI84WksmFLM94QbgXbpKN8fVB3zC/Z8x0Vx9hGu36XX85R2b1+9XL7frZZPvP8x9vRyRHbLD/V3vLu97b167vNLdxnZ/VVSM3ngwHRad/yVqJZnfOJRHUOak4mh2O9bMWPyb/uRyfhTUCTKOsff2Dm8zem61K++28ft26esk4X/SFFHeqMq+uvE4gbM/53hLXVOX3lotc9lH9rc/OrnFP2/o9+4Gd/+nOf/vivOpuZc1lYtCi7BOM0gnEZCLx6EBgE2atnLsdIBgIDgYHAQGAgMBAYCLymEIBKMlpuB4d7JP8c7hDKXecA+YcMIInjSAAjvCedY8Zp3kZ1Bna5diKFwNNQNqfvSIIgYCxvXZc/I5Nm+RwtA1EzfyyG8uokaiTwJJQkCjUo7UVZiQylu22qwgsty/T7VfZI9aDdvkatZr1JQJyxH9JsJgNcZWyvM8b0o0psaWBRiphwLFUmQmB6jnoxJAju5FTpNiNpOouLYL/GiQ7TgQyY6W/2Ur7mhy8htKjTJwcnvCE78DWFfraZcfPtr32jnR0eeSgSwM+KfCqpZM14uyJxRjlnvJkMH9QlMYKdtGqrEy/JjAF3MuJCZsXHjvukyzGj98xD22fgEB+dbwgbyC714uTFVZvBBnsydI5z6v/WN38f4mZuoY+2/h+SqYKjeFlszx3++R9PldJOZmEiUWQfVszWojjPlkW/PBWGkpySbY5ZsiTrg26SISZ0FdTT2qPLKdlfm3zMgK1ypQVCZ77HlsqbL7TDW2SOcd7Y5vp529lZbdubq9wzPyLLYfzZ+gkr0130kHfHqCFQiG2VrjkW5wrBEC8hA4toYn8sktM7Ba6OKePyXm2ZgvLNr7k6q+R7IhN04rPT4XrEQk3NREhmumk0o89z3ujEf/PWFy48i0/6ct8zR7WhDxavElcW3wN1Bn/1se42on+lvfOdb2tPfvVb7ctfe7Z946kn2zPf/Fp787VHWEd2uiD77BsiD73OumeZSRw7N2focyyzKWOznw1Y5CkNOmDBdsfIrEHPCHMcfhhAcmx9tebdOc376pZM1oNnCKY7iyDy9Mkp+6qkTr82NiQEI9bWstVygcOa88vfr/Ptra3n19fXfmlrbf39V69c+rToO1cMSM4gi7STk6Vp/DsQePUhUG/Tq29cY0QDgYHAQGAgMBAYCAwEBgKvbgSM8BLlua2MMPoqweF16vL/3xJoEh8bvX9nMQjtP1sNKheBqQEl7SlT4NllDDaVNfCuUs/TwyI4VW75ZwDazzfqAWzXubDVNdK3B/Zdtvv2oGy326/atCzLdR3L14LoIgywzT69X13v19Xbu+z9dsCMIB80goFty77YN+ckQbq88ILnj9EOJiGzxBr76rVIRpmBlvuOszLee7Uom3v7VlXquI3vU3sy2SRcJiKky+TsLGT6mELwhcToykpndBWdhf3wA5AWq+3qlcv5mqXESy+Ot2fspA7/OlZegwfEhtt2ez+3vEn/qCUE1KRM+Wz/zBgvbGTdTazVwndk1F34FUFr5pIEidolV1bIfjpmS+Xe899u957/Zju/d7PtnHGWGhzlLr9tyLF1vlrptsrIM/UhSPHVJeWZWo4tNNbSuPQB6jm+znPWG/MxtTsUeZ/+M9tNPwvTaaBcOkalS/wv1mV/D/pYL3pN80yFMrVts9eBKD7U1ywlq/CaZ2W8WrpNx6R/wU7yE13KOGa5TOfgyqWd9pY3v5FHtiNCKj7xuc8yfWDKOnWLottj9Tnzq3Iwt7vEmD/1SVx33UqUP0Vy+9zbrNeX+37st/Rvh+eH6a9/SzbJ/PK+P/vemQ2mnHX6Uu0+r6ePdkovc5n1sXaCrtPt7W12X66tbG9t3NzYmH2Uw/nf9+ILz336b//tvzX3/aSYeOgg+X33v6cKjTIQeLUgcPEX6NUyojGOgcBAYCAwEBgIDAQGAgOB1wIC0gthD2ZrG1tn8/OHyZu4YmBskXgISWAAPwWdBuk5nH0JHduWi0GqxXoDV6+9zuv99xV8m1EGHxFZ+yrTA+YKWNVFtgcBZ3xRv4KUPE8+9EDZOkuyNyYZn2YGrDXktKvTn6V8g+CYsnl8rq2Vy/4XYouzvewIyVN9jeaxO5E23srF+Ot+KW5RHrzrATqA44xyoP5UEY4j2yF7hVlwGXtr337m2dTmC4cE6skim8ZbDfzLsxgY+Cfj6wGCy1Ad9sJ/cKbk+bfu81j4uQq8i+3uLvgVNrUu7EYKjv+gqoTMETSbT4YjcyHm+ODZXZevXGo7u1vouMDdjLee9aZ88FQvOPlVwY6vfVwP1XRhP7Bj/1Tf6E8WJJ4zuvv4CMYCidd1FeFT8919MdORRCC/QAjh5VrBBlsq53fvtr1nn2l3vv31trp/q13ZPG/Xr2y2HbZUbpLptE7qm4f2z7DrOvbeNV38yDTf2VJYZF1/LzynTn/yDHSMFJ/N3Jswxr4kESxSfufogAENLs5LxufcUlVfdCxb4mNhOBQVFMlUuBbZdP+aFBeF6zw4e0lu5VdK0l6kXxFlztMxfnX/HW/3R93+XJtmk73j7d/X3v32N7ezk732lS9+vj399afyXpwen4SIOz6Zc64ZPkrGUtTpe9Oz4WID/07AppOMrsnghh/6knVG36qr9ViH75u8JQE3q8P08x4xN+iXNJMw29jazNqYzhTThejz8H3JMHVrz/lx/WVs+LqxPiNJc8VtlZJrX4b8/Uenx0cf/B//h//2xV/86C/oP53XXOgsy0xGdI9/BgKvZgT8vyyjDAQGAgOBgcBAYCAwEBgIDAReKQgQqyVYMxo1eFu5euXK9dPj+Q0Cv91kA1HZiYge2BmkWvo1D/+Mz+rqeu/rbzS8VLpNr92e/XzuPwPWXrrMcr/eVlcC7hrz4mp9r1vu7309Twd7I9fb7ROyCF0hgNiel22ck64up17vl6/2679+BpukxLIP9uk6tGUgfr8evmB56xYHKm0U2RPyo/xLX0mJqfR+KNBpB8vPtJ77A3XtJ9OFQN/St8N6L+FRei+yh0J62MavE2LBZCKuun77Wd+vcRWC49pDV9oOhMQZB8FLmnU/Ow7a7XUPjj9E2EQqLctLgPT1YZ/eFkLXeZh0SnhNHEx867a82keY8DjkzPzkuK2SObbPlxdfevobbf/5Z9rsdL9d3lxpV3c3G0eONY4ey965c4iiEGMYSgYZuiRe1Fl+1frufi1fQzjjV/fBtow/5CTzCSHmnGR2wEtiZyFDfe9X5JXzX5j2rCvxKBlnqwhpnyW0tNOzx3q/yINx91EZf1V852pO1e/XOaGp4lPHXVmJ6HwFFWmfL13eae/mLLJL25vt4N6t9slf/qV2engAVpVFJinvl2zD9WHKPuo7p85737EQZqarTTqt18fITfI+u+Yk0ZZLr7dO0svn++fn4n3ta9Z5WyIEz/HRMxnnzO/pxua6H3NYR8/65mxtD47042sr5+/D4Q/8yJ/6k1//u//rj7uI+HKGg5l7Rhm7Re/3adm/cT8QeDUhICU9ykBgIDAQGAgMBAYCA4GBwEDgFYMAwZqRZg/ZNo4OT64SoHI4/9rGOWcoZXuVMTnRuwGj0anZNx71ZHXfVmUAabBpCJ7rFIyvot7dmRxdhhUaUeHX59TlVVk1WXKfeggVyQmImgTpNqLHQL4HvD0otmsCcmUonlVkm/q7H179VWBa/kDzIJOBpZ9BsHoM8i0Fi3cSAZNvPqG39GgHcgH7/Rykqo84vtdVdTlvq+tAvsv1a/yUn0QfXhcO0at/FxhknNS7/ctZu3n7DrIE704CjtQYixSJczrIfPmVwNgCg+BeQ3Q0tBcB4nj1Ewamftzn3Cek7Ot/1ClBw11kKgsLxKRW9UE76NbG3M8HSnopS1mbssg8kD9fwzw5bG947NFkaJ15YD/lYp4kb8pntNa8oNMiseOce8j9Ym0IsnNsgzKQKR6Kn3snQp/xL76LCaWfOZexMfZT/FLf2akzMG/r+K9J0M95Yreefa7dee7pdsaWyu3z4/YQeyovcxL/9gZWGXTWjYOfBjxZR4d+strAdXnrp5llsTetrzjFP+Wj52QV6cMkBJdscZ2ElKG301EZY46Phz7HeUf1hWKd8qJXrlV9kUycO0a9NemPh2cyU64JhGMH+9E7yehPyvRuKheMfOZ9NtNL+cwFykNogat20B6S8M1vfUt769O322ee+Eb7/Kc/2b7vXe9tb3jn74zdY8/U2+LWMbl2yczzfDOfteRZfW4dltRCISUOcMZeZRM6F9qXZLOP77jvSl8r8W3C1DqzyeoLtDVmZUNkojZrDJ813bM40beyNlsn4c83xkwy/01248n62uyz6P8H0KE/8xf/wn/x5Pt+6ifxMQesFeh6i2+FuL6PMhB4dSNQf7Vf3WMcoxsIDAQGAgOBgcBAYCAwEHj1IFBR58V4Ni5duuTZYxzQf0ZoWsEihAex5kUQ3oNN2w34Kujz6bs/974lUQSKdV1eQsXnB+W+m53er8t3nct+eG/fXrfsn/Jdx/J9t/VgW+/b67vObter5KClyyzfW7dcb9tFhk/hZXuIMWJn9UuO9KC+27cf7MACI0TaSy+9lDrx68RFbNGYrzBaD3Gw7EP0eRg9bR13Vaef8jUt9IOAkDCqoUGKVsaZ/Z06+5YuHEFOOxaJHKxj/yJ3wKy0+uhB+XLGofccfd+uP3w1RIz9xL/Pmc/LRd86DvGTxov5qvW3aMedLm9d/6WOfl4lfpbrY0vSZOor6cEKqmyo46N274UX20vPfKMd336hbXDe2KWtlfYQ5NjOphhB8koMQYKp157J7HJbos/T1Tp/2u0ZXQ/6qR4Py+9jU1afMrcSXpI/+CURZeljyEPVpF15twvnDDp0WJSV+Kp7t1YWKUlDfO9+eu2lz4l+PliiDztkS+Fj4VxrUELp4v2TPPMnsWkWomM3c+ttb31Tu0I22cr8uH3ilz7WDjjXTfLUcnR0FH8lf08guk4gyLhQ6u+Ed6cntV68X8axP3ef3arprz/nXUFI//u9j7T7VUkByg+SLBPLnMr6zZEl+0vgJdV4Oygcwm+C3OlsffVpbj/A/27wE/PT45/64R/645/5Oz/+t/fZR9z5AfsV+FGvl6MMBF79CFz8X4FX/1jHCAcCA4GBwEBgIDAQGAgMBF75CCxFvsZyq+t7h0fXNk9PrvFABlkFluen7gwiPCSorGwLg1KCYoQkBIgvlwJO740FL1RXwK9+SYMpoE24WISP7aivrCuCaIvZS9ZZcu2Bu/X8yoaN+kEsS/Csnvg09dPffJkPsQT0uXbfJEmsr6A7svTr12RmKRCNhrdk29BuxknVTfEuT/E9srQQMVs6AaG+NSJneIHJXo2rqJQiICXELBe2Gbd1EGK9SDrZR11mkKlv7x5b08yo6f2tlKfCz2QCcWsGU9onciT6zKqhT+ozLWW/7F3Y9MyoTOM0Jo061sxNzKBDvfo5zRsHheF7rFBPdg57ziRF1tb5qiiZYjZ5nt0qexLf+IbHIT/qS49mr0lYJGMRdtAhJcsL/c5wSC3VkgmW/+BarasH1gkds16Uiq/TGqZ+Df3a145rSCNmIq1z8NsJ96ecMeaZY6se0I4PJwf77d7tm+3ec8+0dnCHE9YP2y7bKq/s2gefPExf8gdVUCUhgDwnrYrjsVnyrHzgjvXI+VeL9ELaHR8KXN6Oq69761ja8XdSWOOivs8dzTVG9aub8WprkZnpvKhDByV2mKrYUmGw0CP/Q71fJKUEu/SRF0IndXPmrTCNSNmf5vt06ldvHu30DRnKeo3e6HRNFDkWjYz5kRtX2tve/Pp258ln2pNf/kL71U9/or3zd/3etnn5at6hmdmH9HGuzOTyT0rxV2AtflEpXWi96mtt9ve5PLVtwqUYNmcrbxIAAL1ZfW4Znq8kKxODasTmOYftx756eJdZ5v638PHmHN6Md+tkY3P2Vfz5yDpfq+TMuI/96R/5oW/89D/4iRNIYf8yCYEa6rK4To/jMhB4lSMwCLJX+QSP4Q0EBgIDgYHAQGAgMBB4FSJAeGkkT+GE/hs3blzjgPPrJ/P5usHpMYdnExxbIuLVMNKfkWmvT2hJcG6E7H2v96qeNBkymxpF6Xq8jzwu9K2Ky31jRyFK15ugGb0G4pbSlRuFFnW5mf6xr/2M+CUifO7E3LJcGAEqut3yJUHzwufyQ8wq8M3z1LHaHKMZVvg32VkQerRIagUK2jJmweEnCSRBoo5sSf0OPyAfaPPrjZxx3w4OjuLTXHP0tQQL2nOlSl1FmtBI/QR/6vVN0ivZX1P/bH90WDyzlww3S686/AZfiD+3DZLts7JChXtteXY8AFw2gm9hUySW1TyHTEMUsmID8u3Spa3UZ33Q1uej5lMcSgeaMx6vlswJAynyo+Yh42Q85W3JddImeuOT66/mHS059F+yQ3JKEijZYM4pmJzO+VrlvTvt8IXn2nz/TttuRxzIv9KuX95qOxszZzf+SWI5nWzIrG2d6JcA9Py+fPQhxA3+IOecnqJ7MT6r+XKjWVtuQ64z/3hfqNdnKdHl4hiXMXIMlujTHzHG/+DDnfIxPN3ncVqzlcVXfe1Dp8irv5NNdJt0eFf36l7Wr41sT2auun9dtuyrGt/wNcvk1IwubJEp9/rHH2lff+FOu3vzsH3mk59o11/3pnZjc6etcWC+h+SrdwbBqt9sW+Tbl3w0QbwhJ/3gROy6tReayzWkvY6Y96kTeEowUtFUfA5hyTXr78wEMgqkoiRnCEuUnTIuP5yhTN5paEak7jKA5xjXk0z1Z2j6wPnpyS/+8T/+g8+/76fZVgmPfZ4vb2RCJosXa7n7MK4DgVc7AoMge7XP8BjfQGAgMBAYCAwEBgIDgVcXAoaHRrwEl2wbu37D/3/2IYLkKwSB634J0AIRtTJjy5zb9iSlKvAkYLY9JApCRJSGnyshLirYti/RJP/SQnxpfLrKP3NIAXVgww65el8BrrSAwWuRS4alCXbR4X/OFqRJBer00kxkcjPdR/fSfXzGtvWOqmf69HqD7SLceojdtV0Etv1csviJnovsrSKerDc6toTsSHZaEQdmWhW54c7VCZNI8oQuUM243bJGBcAxWn8LGbvVQe/r65vt3t5xu/nSrRq34zJbyH4WyQLmRrIrvqqS6mS3OWc+oDtlFX/SD6S5kiiz0JX5JfMrc6OwfbAVroDHtMt6mEXklkrPr1orGeU0hDTyRWjYHkKKMW5trLcb16+yFtiaSLdaamAAoSROizUWPWVaP8yIk3BRxnFIFqaeNsdqBpGgeV9rrK9Z1w4ZY5NcfPMZfXyUoh0e7LXtrY38jo7utW1ImNN7t9vRnRfbDrvtruystqvbM7ZXbkB0od8PC2DHJLueVen6EVr9sfiv68BnM+Mscqb6bEJTMumcK0ky/RItnuch1VwTNbaMF4wjg9LK4FN7vUOSaxhi3lLcxtEAACAASURBVLgwJlc4iWshXCXvgpVrSb+cA20hn8xL6+jhXJrZxhH5aUeVw7v40S6BS0dquUzPZ7z//p2Q6M22zswlMihwTZ5PmWD2Yfbwy/lltaNrc32tXbv6UHv+3rzdvnmzfeYTn2z/0uVr7dJV1gUAbW/jj39vJBw5yqvw0gd+DOwi8xKs0Ok77GgcW0hHvVfW8XnPrX9/qOSnnP9CvOXDCvVxB7ZKhikFI+BakcjlNUIvsmQbHqH7Jp2+zFlnn2SufmVre/MLm7PVr//hH/hDd973M38/fyPRy3/7C6YNQBllIPAaRGAQZK/BSR9DHggMBAYCA4GBwEBgIPAKR4DdZhVwvv1d717f3d29enzngIP65+sJtgkSCRTdjXROrJ1SRA8VkjJGg9bm1uA88iXIv+qwGGz6S5YUAbWl9NfVe39rbEFT/wzmofft13Sa/ul1Eg/q7QfRSzNZbO82+3Ov68+297F04o+eC7+Ui+5pDL2/dZbeN2wA/aoeXyJfRNya/GO4nPpaHokqmLB/4dJ11nMRDdUfrZAl2rBEd/yt+729/XZQ2X2QAdIZVeIvpIIleiQo0JF7zK6sccA/uThhUNAX+er6wL8Kd18dIeMi0M8HB9Qv8wLxhQbqy37pAj99llSYSBkzwbodx0RaTtvi/K4dMoX6+K33XlSUlUniX8gRstioV2Xag23HWrKsCFsa478yFnVczE+q8o912qp2SDDXD13mYLnKuI7u3Mb0EevvLGeOPbS12nYZ6uWttba1Tj8J2vwkbiRkxNC1ICaMk/9IWPXxVBuEmNtL8a2PRWfIh8rHAfzYgfgGI3RLZF1gZp9aAxkPssHH/mBUw7XOZ7XWXEtYSayZrSeOCmjb+2WMUkc/M6bcNpg2AcGjLmd3tzVqH+0L/GyXrOs4d/nMMeveesuFv/3eNohR3vVT1ufqbKNtre20p7/5rfbkl55o73jve/ja5UOcRXYCSbapY7zfYtzaiRloXN0aSwOQ13y69dgPAniYfm3FnMY7jVs/4p8YTHX4eZ4Pjpxlr+weRNxLyNxkum+BHF8LaKcb7BEGx/PVtVVfqn2WznOM60ubWxufubK7/vmvfe3pOz/yp364/ew//hlNrLO9Fblp4NYMciwojH9emwgMguy1Oe9j1AOBgcBAYCAwEBgIDAReqQgYL/tVtvav/5v/VvuLf/mvzMjYuDKfn1yZnxzDTBhwEnHCapnF4blWkh494PXKf8nkKAIkICRIv4Cjyxqc5l51ScGZgmXkU48t/yNbUe08LfXxrCMD7wsiywB46usgJCV0xhH57H1KBfAG0Gm2WuKGizJdrs7qYhxmvaiY4rVs1L1fxJMIqT6Op0iDi+eyGT5D8ig+lK6YJW5WJyH9Qr83ZhQZ7PdtdnbrmXLdP5QtCEmOB2+3OBvLg8rDVUnMsA9MzcmgAicJMLZ5cUW3g3DeqF7jbCVJCcmckFDq1WHwsWjPX3mditSb+WPqlHNgVmBkYC1CrqI/JJ066xA07Hk+V2X9nJ2BPUSUOiVNZszxpa1NSLJ13DiIfpeZ8y0LEZkQIGgICRcRbImptso75cQ1hBy++Cy05Vs/hH6idfHNWY+/kw2/jqjOUw6KZ723o312zqH7dP8W57yttN123K7uQOSR6bRFZtxMX0wBA2e1Ss444hVT4HAk2GEj9mmrrDHniDUDxtrKGgYLXT1bOW1rmxu0OWb0gqvt0cNkZYsu46EbJd5DZE0kVrDo81TrVL/Ew6vy2vA+M5vMurIvysnsco2oRzHnHDvOAV3plc40OJ5pjTpGquOvchRf5diym7oUprBC8q+oOy9rELM1RrbnUnd8ct7uHhy3A9bw+vYu6/JSu3vc2lNfeaJt715qb333u9s62BxzLtwG68QMVi2e4rMZe0KetUhdyMR5fXWUx5TuC2jmuf+NkuDFR1UxVO7Pz475YunzEG5Poe9Lm7P1pyADn+b5NlNxSO/z1Zn7iM9O+Lu0R8e7G+trt//W3/yx2z/21//a/tNf/xoSgpKBTxOhc/YUlPJn/DsQeC0iMAiy1+KsjzEPBAYCA4GBwEBgIDAQeMUiIKki6XTe/tgP/mB77A1v3Pz6V795hSD0MvEe5+gQ+RH3EThWlMk4CalzHlAfssGvoXsPjA06e+lBqm29vsv1LJsu2+t99t7/oJUngk2K25wsbonTokG/LZJU382OsgbQ+ma2icG5zxJFvSzb7P51XcrYXvVakxjpcXBu+ad8i7+46pbL4AFcdE1fnw3SYxtsxFp56w3Tk0w2qStb+ldwd5/Mcol8thdyLtPaRrt9+3bOaco5YPQo2e4vGiRaGGs81BkZBfRK1iCss3kWS5xLnQfIW9xmWayKYurEf7Ol2I5pxpD9Uy8JRoZXvnAZbRcHm0dR/EZcDGKv5sQ5uLLLWVOuHUknbdChjzfzho1gRotj57+TnJllhUfkIX7KR7kJfui234r1EmlxFx0c1OYyZq9wXLOPLomHJIwE2cnBPa6HbWO+37bIatrhiLUdlt0G/Mg2W00lHc/cjheyVUyoim+19bXWg+eMHeOhWPC2QOx6lQR1HZ4cHceeMG6QQXd6crRY2/qEVPSeQyq6QIrQqbHVOMFM/Gv1Mz7u+Cpox3eezCzfCdcd46ZtRXIJ+9GfL4hK2pnBhZeCMGHf8VeuE9HBNHMxzS3ijtklmjXJNX6Bu9dlXT73n/p8a0+RY0drO2J8L907bIcQW5uXHmqnK9tgDjkJPl/7J0+2h27caA/zc1ul55FJ/cVfrpJd/NVCt+PUfsxOtn1PtVv+glzhVX/C3DYpMcbrkXVzxpq4xe0XGc1HyBb7+Pz08GtPfOWfPL+zuXUHRYePPfbY+dHxwXwVkvTpp7/ZvvrVr7Yf//H/pf3yhz9I87nwkYaGQ5V+5/bM+BHH6m78OxB4zSIwCLLX7NSPgQ8EBgIDgYHAQGAgMBB4BSMwBZjHpydbxycnV4jpL7GTyQCUpLGzZFpATEXKIN8ScserQbAVEhNGqhOXZn0CadtSKlA1wykBPnLSN6s9kDXop08PyL2PYvRaur4iPwx7JQYkH9gwCOlUHJ4heBXrK5CfAmRJH2NX9KorZAlXZUpnBbZmR0kuZPMc95ZkLRGMFyFQ/dVvEZVkakEU2e65SOq2XTshqhB1GHZJ1hlkAVE15JDnTWFLOxBQ8deA3gwvSnybvqZnX7O4NjYgyNh1dvulO2wLhAzwa4p+KRL5wtI7CgbpkvFquMgv9OpIssdsk3R0jP76vDC/RR6kf8ZpM0V/kq2FjjOyoPg0ZcbYx1qYTOOGYOpf8pQsmrOtM3Po2Bnf5Us7bYOvRc5WOXqdbKKsN/xQRj3OSWxmOB6AH64WJ/DTOucTecm7fhYVg4yPzpfn5SkjvhbJQkvXbb0qJG5Ojw7bC88+3U43V9v3PXK1PcR2ykvY2wHXTYjFGXitQHqlr1+rdF75TzKiohOHMFO+I8saDzGFTbPITvmgQdYGJNzx3lHb29trOzs7mf/VZEZNJK6Im+nGpXSLAz6Cu7r5p3xg2rJGpuecP1fDrPcSfOMLvnnNeX7gEUQdN+2uObQJyaIomznWgalAJaEkw5uk8UniE9zEg1cvNmbTmo/f1Mc+fp/48QOKH3yQHCNhrO0x3y/snbZb5Get7DzUVjevtPXVzbZ5bNbdWbt792574vNfbCvv/R3txiOP0Jt3i1HMWOu+M/mqZXziOfOKP/zHNRMajnFkZXPNV1aRdRD45F8MMUoNPp+szlafpd+n+bv2oYPDvU/9kT/0B+987tOfmrP989TxbW9v0xc8IVv37t1DjQPmBzvqCmN35vSi5VMZS8Bpc5SBwGsbgUGQvbbnf4x+IDAQGAgMBAYCA4GBwCsWga0tvig4bzsExA8RGHrwj8EykSFcA4FmL6nKcwXrtNLPgLsIli5nH3/KW7w34PTX9YUEmQJs5XxWtTK9T26mf0o+HaipjJLs5ONpWa/iy8/eS5h0n2y3LMt0nzzHyOw2E9aqXRwufO79Fn0Zv8xBtsNN9Jxt/iQkMm4xuICwyB/JGzp2PWZmRR5d/VynjBcdwQYiRXCsg1cKiXAO+bLKVsCuI1fIixyDpKOW7p9EAhNssE+H8kvHBZwikacHnn9lu1ezcKyXeLKof7qJTPV1fumnfvume43L+thTAj1nHkavAmiKK5cvZctiHid/bMNq7PR1Y3svsT+5kHbJVTtZlxtdcP7k7upg/I7Nmh8jUAxbbtOrsUDwnB61o727bX5wt21ubrddzmg3a2wTPRuQVX5zwC8oejZeMpbUEU2lq+Yoo7IihNtKcK55Oz4+qvO9IJQOyYS69eLNZJDNYFY53qqt8yXQNSY0fqLXLY4Svx07D5/XhjxfX79FQvWB26dsZa3RPwUQknXJo19iNBPLLz/yFlQ7o+iiVngvpuqwePXw/cwbsv39/v/Ye7cY3bbsvmt+t7rvXXufs/e537rbbXe6E2KCEzuAcEBKeHAEgg6WUBJw4hBIFBMJRUJIeeAtkRDiAYIQICGSt4BAEXIULm+EBCNHDggc28fdx30797NvVbuqvvouxe83xhpffXu7T18cd/eRPOc+61trzcuYY/znXOUef485p/k1NjVXfE8caBjzILEJskrdmT8LiM0FuxieM073L+btGx+dtfuXAn0EdcpedOtpm0H+ziDBLtgP7vGjx+1rv/G1NuVAiuPbN9ue+5VBnrn0NcaQuX+FPO1Co+ijot7UZwohVymwxawcczg2wLcVOp8SNfYVRu2XHz249yv/3l/8uQ/+v//7H/gHj4m1cFBW52eXOfkDEv6fBXy1wAEfl1SxFlc//d4R6Ag8icD1V/hkfn/rCHQEOgIdgY5AR6Aj0BHoCHwSEdCbDo/afaLm54uj6Wj3aL6+wBnVSadsTDyM5AaP/tMZD0eTPNO2U+27dS0fnNGNw41/OTxnmc61LuZ0kBMcjMLTcd048isc6pIZBIC0Unj21wSTPrn7WoUpQWTY15NRNBJFUUPyxLAvayMnoreUhz4mrarlnPq+Ftm/znf0PxAxBAkFkWXUXGFyNSx10/lm07YNkWCglqccBPGFQMkO29dyQPt1P6tK9hOYSzxQ0T2XYmkjctVNnc7P3UNcDO1NWUa5SB7wLrs3RPhc++9l42B7Kl1dxj3xVRh1QUJ8srZZ5MUlVIllRWVFYyLdIt/IMttZx/qkIFAGQZIZsFLt+HAPuygEDKOo3GxfG12CWn2LgRFVMccgQ7w7QKGXuGNDaZgaKQ/xyLwkui4j/yRRjAdMXeLEQp4VLWYnDz5sDz98p91mJ/67t/baPvuC7aPXHljucrHfVOh5hc4RDUgEGdnIGwcJI3FkP2tOtcxoNCLNkOuywJi3kDqEIsX7owcP2Hsr840ic4+tMNH2tIG44XvQPpdFOs5JjgFM6j/gSQHznW+SNrmM1HmsjFx+Cgpox/cRczaJ1zWhW4hGlPdr3ATMsZL60VDnzwZf4aQvh8lvzDLbm+dlijHh7rvP/p3wv9pPb813EJFjjN/lFXvnXazbeyer9u4ZxN3kCFLsGCJywob8EIl8u9OdadvdOwq+88G9++1rX/kqz6+127chzxgLP7+IwozesZeMMYcn0HWMg3oYSantPk8r4i/VjVbqOXHJ7GR8bzqevcU39JU/+zM/8/Af/tIvKCT6YG1soKRpMY5hL3g7EsNzCOs/HYGOwMci0Amyj4WmF3QEOgIdgY5AR6Aj0BHoCHzyENDtZQ0ZJMzzz724wwlxx/ibR+opqYAjyeltW0QPziPeYTjCOtWRwmHFcR6Wdel8bsqyRrzrVJo/tApHdChOMTqm1Cln1OgTyQdTtU3HlAwYCgm8eg8HvyJtkJH10yOO5WchJeXE0rvh3Vv153PoDQDSB+ZX5Nh2/2V29V32xt5o2L6dL8GBOsjlJ+6D/YCQhBdl5BvRVJjZvmQUGZZ6usyM+kSIyX+9/c47Cg4sQtagmKRVnORno62k/JKbSlE4tBnHyZbQJjI/jhD5UV89IRqCtTEPTFA3CKAIi1I+4+4G/273FeRL4KamT6bAiTriuiLs784zxzQDL5bV2auEhul6PBLLQcWN7mWD8rJBEnPaZJl6u3xVXQL00HhLLnXiBEVIlMX5WfuATdZHi8ftmYPdOK1yD51Yadl2AXmH+xRC1iV9buivoi4X9ZuIvrBHgoriCM5z/yyjv1bMTZ8l/mzkPLo4m7cHDx6GyrsQYy7dU0YQmugcuJZuag4xeI1FNBvss6Z4DcTW8L3RlJTfS4wdfYqrP4EZ6ktKO4KWq5PJ5cBGmGUbqkejbBPtopbviXfqnG0dA0YpvlPzN2NCpwwBwsGJZwIHiRKbtpPFBHJs0d57DH139Bwyieqb7TOfp+1o5yBIxAlLuN2bTfvmkImPHp229955lzGYtZvHR4HJmAMl1VdljU6z31zqOY2/W+6v5lJpye8k/CDE8m9JKG5bvq3FzmT8/s509uav/cqvfuUf/uIvXIwJF8QedhSLyciETJuv7RrA6LeOQEfgO0KgE2TfEUy9UkegI9AR6Ah0BDoCHYGOwA8YAd1XncW6WAK1PsbtvE3E1p57OqWDC7UTESNG8eAIQwzYcCZhkB55SKB27tlFabqU19aVk1338NgplhgKJ/e6aji/yq18iSP3O4q2dhwO7xA5w3NEzHA3CkmSxr5zLzLrSthcsYRNJzn84pDLWxRWH9Wf4rOeESjVB8wHUp90kAfiBlIxCIxB/kpCgnaqk2mI/lECDrxLs2LJIk9iCw8TTrx9BhFGJJh7RcXeaJSZL92Re6KlRPub7exBHECQvQ1BJt0BkSJhWPZ4N4IpCA2e432wP6UIjSgkJuapn8RE9GUG+sX4QyK5d1nVVK5MWPB9EEbuSx7skDCZwCAikTBuBCGCEnFJrK1ZNnfFBvJLyLEDTrC8e+dW7EwW0VfIDf1prz2SWxIagZt9ksTDOmuYkBynHFfbRxkKexKpc8J2MQ+QIUESZNIQjUVAJKghBxDvvf1ee/DO19tNgD5i6d4++46xbT5zhgw3RUPeKCLXjOiS2BMnCSFNddzUcUlU2JLN/Ykg41n97H9BBJtEzYioMN/PLy7b2ePLINRczjxlWWXYjG3qd8VebEYK1r5uHpQQc4r5V0RZzAknBRjFkDowhiJuRojHSOKeJJJLNhO71ENKS3mcVhuHBpxL5PGeifvwGLpdT+bNfBE9JMZYO5+nXMqXDLaNOC3kl8DukvFcULaa7LXHF5P2jXvn7e1HfJO3X24v3XquzSFHT8/Po38j4sRLvU0zyMUp0YhrwD45edzeffe9IPJu3TwCz1nbJdKMGcHm/vTNRv/qrWYRIcjfKccnPkXuktdBUiPXb9vvbTadLiEq7+3vz946Oz/5GgN+yfzOta68UNWvVENV54mknfF9IFsoeuoIdAS+OQKdIPvmuPTcjkBHoCPQEegIdAQ6Ah2BTyQC0jSk0WR2fPP2s4tVuwMptRuEy1CSBBlusSQHjv4MNzSW8vFcDn6ZpqMcjungWKfDHG5qVdncrWuqKK2SFc7nUBYRS8NzOvmSYqlYEVslp9q5vE5d7bVk2o/PcdGt6m23i7bILaKg+vJehFvU4b3K1NtnrQi5dkKq8nquu3XS2R7wwLF3m28XcqmttEDuPyUBZV4m7bUtZyVAqnDCIYSV0TIffPDBUMMbhIn1bJXrFqPM5Z8RSRV6k6Xtgw3h4avTQIIFLUHZyKVnyLmiE6PVYi7YVPJmSBJdGXWm/fYriUjVmCO0C1tpYyY1vHu4g6c7KnNvutfu3LpJH5zgSI2wPXTBEnQwFY4e6iAhlBgobxhHbUNu1bM8CBZqqEeQjsiCLot6ammdOMiATfMf37vX3v71X2tTdDritMpbu9O2Bxy77As25bOYTWfoJmDRkjmPTNorV1wRRk/Zv9Fv6uI+ZRI0o9EMQuikXULCuWxSru3sdN7O2c89lglyCumK8VzIsnAtIRsliOhEuEJWLLGkD5cQSrql/aItPuZz28wS1VGfxE0aO0aGORpna0SZ8q0A3lzOIwloiSxeok8LU26IChJcLMVY2yvKz1L1sG59M8SahnxJRBFbsmf9BaFj7ILf4AXbfVYEP1hN2yURYwf7t9rO4XE7uL3b9s/O49ACJe6O9zh4YgFu54mz5CI6Y0YswXz//fcZEzJuHrZZ7DGGlZoAjyX+qyVfEmNZ5FgcMKDJ8vyoiymJBCLA+4LXe7R674zB8dvyRNHsTQslx755UlhPHYGOwLdHoBNk3x6jXqMj0BHoCHQEOgIdgY5AR+AHj4CusheuO7fRaPfs7OzOePfoDlE4uJiSD+H0D/W8wb1IDuCw6yDGHkhkB0kRIrIOrvuGtLCNdcuJDsdycOQrL+qHI5/kgK59EBA2JhXhlpFCSZSkg2o/tEbeBOdcJzoiuHTPjSgjP0mDJBfC8dexhUDyn4ke4wkOJOqbJyS2Kx9Y+0z2lbVxysOmjJwRQYXEssahT8slOEy1j5TkgnLdU03yQhtr2VpgSD/ZgzQX+OP5pxwia7AHK+MaQ9ycsIfTPQgek22iHlFk3uNETfKS2KBPy10eGE/80q8pNlgXAZdVSoTp86tTVBUn7aNMvWAWeIl24kNh9hV2Zr9G+lWStND8IDgH/GIZqTIvIaSO2Qz/gD3Irogqiw5Tr+Vgc9ihbr4jVETMM9W9xiXGUrujU9VFX3SxnrY6ttmGPF4Us2D/r9/45f+3nbz/jXbAnmM32dvqxu6kHTLzCUyCzNM+5j+ElVaJpRBIDI/RV3nWcd+s6ENiC6JpAcNs5Nfp6Xk7m6/bw4dnEfF3+viMPePO28WcUxEB5t7JHNk77cjjSOlbpZawVtBBnPBJP8jWcGUbFWd/cdql0Xt8l36Hfp/uP5fjTD5laafjIVI5/2reOeyWuxeekYrOJskn56mzy1E1uS9ezBFkpBwJNV4AIOYuuFgu6RljgL6RriCYYiyxBQwuiP66ILLrhL0NV5xSOb59ux2ydvXDdx61+RJykBit2f6sHd6YtIOj/XZxcQHBRRQeWLrEMglo+nAKAoYE1ppGH3zwYUzBCX3s7nEKKutgl44zYx768LeAJoFL4RfRr8ilnP9XAH/DxqAwXj1eLJcPDyY3H3/04CPIMU9Z5SvG/DSoEMk3MwNWX594yfL+2xHoCPxmBDpB9psx6TkdgY5AR6Aj0BHoCHQEOgKfPAQGJ1DFcO4n072jo6MXT+frF3Ai93QswwkmfKcccGvqgMZWTEO5eTrrEjjpnJuT9WynjHBayUtnFZJicMAH+VG/6nnnv+r7CZnh3Fuod4pznBuZW18iQNc1Hfty6u03dC+3lra+G1FlbU8QdAN85RqXs703WdqSukuMmKr/0rvebV0udbZ7sn61jb4lb6ge2qKP0TaSepUCM/Dx5ELJGF10tVWu9kpmjYicOXl01i5OH8PkHFIBacGFaD+YUyfrF8EWgGanyMsyWQCWqAmnGLgkDrlhWwyAAtHLpgAQkTgqLRgCHHVknhxP7lQXb9tHOXUics139E/ck1SR9Do6IIqIfbhGS/bscqmm9tHeuykx4hl2JJaQkldEj0rVGFi32tgy5ha6hJrgIrlkdFEkbleXS5Y+ztvX3vw1lld+vc2IGOKsACLIZmzKT/QYdafo7Ib3E3A06s1N3tXfS0lhC7rGPmbkebJiLOMcSJ/5ckLE1KjdO71sp3NkgOv64HabHd1l4R7LNyFoFvT1gO/m5II+kTmD/BGqHaLYtG0K2RQRZfaHLvYpsRV6kBf7tmkbdfOgBzO5nDfkSRHld8fYOCRgEYQ2kX8mD5Dw4ACj6UAz/0mUOQYqYh3x4solo4wny2mNxzPFFl3IlHhaYlNEohE1t0THOeMZBNmavwssrTy6+0o7euE1Tq88aGdv32+XX3vUTomuc+muRODx8Y34Ficwk0aPLWeXKVO5XB624VhE5B8KSTR+eO8j2jgvDyKilZmEvtrmHmR+B8NcJMd5E2OmvYTBiQ+HdLB28+qUx5Nf+ge/ePnf/82/mfN8wEcbe+oIdAT+8RHoBNk/PoZdQkegI9AR6Ah0BDoCHYGOwPceAbxg3OvxFG5r3I5vP7O7uFi8sFquX8SH3JsPZIVUgZ63TmUlndaIJMNpT4JHEiNoi6giYVH100nHoUaeeeGc4syaqqzq1t2yJEx8sk2SEpIQlV99rFgeZx3idkK2pEUlnWLr2Z332BtLW8iKaCfkSUDZwXbflEb96hdNQyTi0FnSySZpQ+jDc0aD4YDTGT1wlYNOW0gEG0kuJJlHf0hMOQiN/iQyMipIysJlcSFbvb2o5WmfM/atkrR59OgkyJbJDvWCyaAccmxBzTjVEp3CdvuR0bQzrog84tHnsEFFtMWIKx7VJXQM+7RD+eYpj2LGEVZjIE/ISBii5RM/8muGbiknxoF3TlE0CtDr7rMQRtjhTk/KNSrRfatC50Fd8QbYIHecK3btclfnWi4bHQjATeRa2qBKoa9dLi4DryCMmCvzx2z4/taXWVr5K+3q9FHbhxy7Mdtpu+g0E2U6YVetGEexFq+AQpkoNOFaclql+iyJFovoKxRasZzQQ19XSDlhr7HHayKgDu+03Vv7be/4mXZ469l26+6zbYe9xw6OjiCU0Z2lmEEuXZzT1g39kTmHMUOPFcThJQIX7A9mvSu+ufiGKJPv84AKSSOJvBU2Ordm6CpkoTPyXRJpdJ44Spy6LDaWJdLGSCz7cc6s1ix7Rab7qYm/2Hkpy1TzSFJshe3qXN+uz1jCv3E7uzhl/u1wUiX4Hdxst196DXLsxXbz2RfbAvKsndPj6gHRdafsPcYhBrRd8D1Ndybt6Oig7e7utsnuXrvcu+BAg/N2xWmXE8aGGR36uKfbGCKR2ccJpZftAXLWYHBjtE85Y4GuBvsaQAAAIABJREFUY5bGGsUX+msDmBgJiA0gISbsSBj2TZaT9ejxejV//Kf+5L+x/MbXvhJzi/WwVLz+GxIADD9AdJ2GF2UVPteF/akj0BEoBDpBVkj0e0egI9AR6Ah0BDoCHYGOwCcdAfxi3EqImc/97t+7xwmGz8E83MVx3S0HGOcvvOZtR1AH3KRjGMu0eI5yiaB6pqwcR8tMvm/LMU8Sy1R18yXl+RzRH5BFQQ4MckpG6IjutaTQ+k+UmUEyyuXpZNuyI5emQY5kGNYTeiqvZH4zGVGOC28XkiVhByYZsSMBYbkp7zjsEBIRuUOed1PhwsPmPYbFtgNmRjVVhJsRPu7FVGW2knQSKzKD7AoWRWmDTCoEgaDdYg6fE8RD5Vs19Fdd20A80COZqbsUiFFHYR+y4s7UiMQ7IDuY9m4DfuJpKKY+hM8YQszllRI3t27eoNpAUFKr9PJeEXA2zqix1CHEkieZcy09y6zrOGubUyoxTWLPMvWbn561D7/xjfb2l99s84cP2jGe2wHjcUBE18zIMQkU8QYZSciUpY1GiGWP6uPebEa9mdxbbAHZZMTUnP21Hl+s2hlb+J1C/pxNdoMsOl+x7f9ot+3t3GhrTq5017UxZSMiGEc7EET7kIUB2aodEhUFexU25hb0dDJsXG90lUsQY+knRNWVyxHBVYJszp5d6r0mLzRDP++5fBV7xIS8JSScJCM8EKW8K8elkRB0I+zS5sSOYpJYe3qn44KAiBSTnJMYD8IastQ91iYz9hK7caMd7R+3/eO7bf/2c216cIsIMjDAXjgruFD6Y4wkxpbo/OjhgqWW7tE2ai+8/EI7ProRc3dvdhBLLGfnO41l3yggIYkACDxJYve+s52RZDtG/hF55pi7Ef8KgkySLE/4TKJL/jRsIhSPBKsY0YArTq88+59//n95/I2vfpUwNdFyEL67pNyeOgIdgY9HoBNkH49NL+kIdAQ6Ah2BjkBHoCPQEfhEIIDHmN4gHuGoffFn/nT7S//+X95ZXF7dYqnU8Xx+ifs8eH6s64qleMEApQNdm7wXqSHREUvbvNPMK/KG53Iir/PSYc3lYTimeLdZJhmVDmc45CgZy6gGVQgBCbWrD33djOhCL5zeETpaZsSJSZ9eef4LciXKcaDTQY6IG/dWSjuk+ga9bEFjCSFT9qNM7TcvCRMjbjJlvSIX0v5rDCSbEgM3azeaRTshKRAZ0TdpGP1jD/rEkkuUCb3sTTJCBoC8JG5ae/c9NuiHmHB/pieShkJkEFqDcLGlk6EO3WoM0UvcqReYD41T5yGfvqxSSfU25FhlKkuAI8IK+wZ5FkdbFQvWh3cicuxLUsmosSmnQt40iirIpiHSCSxdymd4mKSO+qROyKEbn2Mj9sAKgkN5jgX5OX5BelAnx8T7kuWU9mv75fm83X/33fbhV7/aHr7/Xuw7tre/0w73J22HTb9mjNFqfhZkz5R8YXNGjIw+ct5QnntUEenGXlVG6Rnh5dLixWrc5pCFjy+J4BsftjPa3JuftAvHeZdDEdmYf8p4nGGf03tHIoc64mFkm7KdQRPIpgV9sR0gdlGODeowAUeXWe4dardDFzPFzwaSjGgpZK5ZXjiKOZsEVJBhEFERUQlGl5cX1Mt357aRYMp2bMSWB4RAtkWUGH1TR7KNEmqhJ3Xc529XnSClpnEd8bzTdvZvtDEnq073DiGodrBnj/3HwIXG7icmb8uRDkgZEUF3EMS04zNnfBqRYm+/+35Eku185jOx7NZv0nmyf8hG/ESVPT47ib3e2hlSkDcF0xGMn5zW4mLe5ry7bFWdJcaC1/UbB/OwA9umADiexMrx+C5G06mz7/GH9z+EgZN9c5ydTvF1aPZ1AnOTqAdW+dp/OwIdge8AgU6QfQcg9SodgY5AR6Aj0BHoCHQEOgKfHAT+2E//NNEfNw8fvf3BszjIt9HMUAv2vYaqgRHCkQ8XMZa34dQHgWMlHXWucKIlIrZSOZLedYajno44qZ43Xugm3+gVHXXkJs8RDmkRIHakrHDik4ZBGm1kM5QxyLGObaovCqJPiTOXlFlNHazjkjmZBvUke9PGsrIonrVzkO+92ttggsx69x6kXAmj/Ol2iqm8JMmi28izfaWqY17u80UEDqQHK//yBEsiaaIbmoT2RB7Bpmhc1lf4kEJGdhzlGA8XRbl17VJcYF9qc3syUqYDMYgJGcoLHIYB8l2ih/2kAnPkuRQx5NqQMsfTMVEmTA1jQOQWSw0pCLJkjU3a6iXhFIt6gyhSMWo5J4ZkjiRiYIO+3p2XpooI9Fldo0/krIm8esieVQ/ffa89ev9dNsG/bHv7LM1jv6+dCbqH0FyiN5N4kRACm4iqQnfHl47CJpfsSbxwOCN55EMIzeV5ltM2nxy00R4nc45Y8shhiC5nXILLFFJoSXThJY32AVucMrIrMZFcNLoO5KIsltdCovmdablja5kb4HuXJHJJqnuSuY+XeLqTWYwnT+MZRBF13ZcrcIJJcp8zD67w4Acj0mKssMkN/03a7Hj4bdVcMTLT9l6BJzY7R2Y79kU/nES6Aosr5hwxb+1yzB5kYLJi77E1z8qSXHRfMknhOWSepOKMvedcIln9GCX2wYfIne63F154rh0e7SYRjGG7Q7TqBHkT1mheArakoMtJtVG1/Sa0x/uY8ZBote+Fc5t+ZyzhRFtJuCvl5VykOQdjTmbTC0h4Dj8VZTHoqSPQEfjtRKATZL+daHZZHYGOQEegI9AR6Ah0BDoC3wMEyhHUQV+3b7z9tfapH/780eVyCUG23gvH0wK8YYgZw3RSB5xdn3VGdW43e3oZsmGJJAKpHF/vkhY6q4NTGuW4zXrkJJe18QAZ4ab0FZCFPx1dlnPuXdIkCAOa6qSvcZKzu7Ql+iY/7oNDb/08iRBjgnCBWKBPI2cGBVI3yAvfy0GWSHPZmPKVpx2VtD3sJp+FZVFe70WMyTtFhBN1bF8ywm4ESXCY57vLCa3ve6XAjzKJE/sTO8ulbiRr4Hfau0TdjCANQm/Ksg16SoDI3gRJVRLJdsyiC+vEf1EYthWhJX6OZZk7qBSb9NuThJCNIWUiVTv6r03+zS97JZIkbfznHJAsc5+tI04efO7ZYyq6VA92SaID0d42CV1kYZQlGRMyeTZVlCFUEYReLWuVUJIskxxN0kQyyT5PHzxo9955p73/ja+0xdkjNuQft2fY82of4gQKi0A8azIXjTpyIaCRUzP3G4vZiZoSWuhh5FeQMPSBsgsUW7Ah/xnXPTbj379zu01v3G6j2UnbkxRiXjHz25hlle5nVuOY+DB7GEs/syl92T+d5LCpB68j9Eq7c0Cccc7RIgyjDnPkEsKr5qj1XU4p7WVEpZAa7WZ+ELmM4do95KgTcwuCMMaGeupnn26cb31PzRRMTnoM+fUdX9CndR009wC7cr0u97XjjSX+mZCsSp0kpBBDvwsoKeitdnBwEBFh05gSMePYa23Z3nv7vTjJ8tVXX26N6XGwt8tUI+rsCqqPPnfB0GWV7kVmCh3I1z73HZtMXCLrPEev6AvCjAi3qE9MrH+LltgTKGIgUXArTstktahc2fbkc44lZtERpZm0LpMzxr8TPXUEOgLfGoFOkH1rfHppR6Aj0BHoCHQEOgIdgY7AJwMBvTt8PFw+PH9O4ruDk/uM74OzTZCLheksuoQr9/UxgiXrcItUhFm+JZlRz0XwDDIje/tZkohD56rPuBshZCq5Ouslp/LDIYe4CFmUl8xtEiKEDD9VrhuM6xvyaomk8iMJRcjKviUAKmV+2i1Bkf1m6aY9cs1XB/WVGKp+N3WCZEp7jXwqG5WUUUWCcS3X9tt1chxaOz05C/lxCiFEjpi5/DOwk+ig3XWfyJSloM4mTzZSW6ELgvfUVHUb+n7C9qBbJE0gsyTHoh11aRiRbTA1SZhIjqh/9h19KRyZ9iOcLq9ky6ggPyRwJHkkAiWhksAr7MkPxa513p4DIhTYqstgm70E7kzboJxov7y4aPdZUvnoo/fZg+xhm8Au3jhkU/4pxFTUgmxhrCTJPP1QEmUGNkZWrSF+7EOMzV+go7YZCWVE2AqC0mWV7z68aI/bHrCwLHDC8sx9lgZeXsW+W9o0g6TZI2Ju/2Avdc7hjefplChAl1Myp2ZEYsW4WS7xJJYkCWOfc25LQmVyLkv2ghwVUM0CsLg08gs9oyFyLJaIXYGH/0ySukaquZyxIs/cR81+iyuKPe8cZpZPhi4OvWNFPQ7sjGR7ToRk6iCX+WM99TESMeaTfVlEfhFxewfsV3axz/gSUAiWCwyUULuCuDxnKewpyy53IMeIuWu7e5BjROKxdX707bjOJ2zuzzJXSW+XHIdsSGH/PlUUmX2NIPh832VjfydfzZ8k1BbjxWI6XV6tZpqg3cqmDiZeY59W9t+OQEfgt4qAX19PHYGOQEegI9AR6Ah0BDoCHYFPKgK6tnrJ+tfhLeNI3lktR8/hrB/GJuA4rDqTa06Gc1NsHVA8yNhUPIzS0SaviCyJDkUZ2ZVESTrE1vW9HM508LOtZeabdJRNblpuv9vkgP2YvGeElo6ybVKOy84kGFJW6hrt1YloJVx1W0Me2M66OO70W5t+Zzuca/uxiTqVQsjwPeQjRb4w3qkYtlhOHpJVEYQkBYjeYZPwyosCsUPsWNtI9qUcqY7szr6VSR9UiQg5xgB1I4UN6gY+RiJJmJxfciQgjWMMbGS0j9SEZIVkA29xGqUSjAEc+vQ1MPUdEsO+qBn9q0Munx1wlOQwqaTTJZSFUPIVoTU2EWFGW4TwH/U0JIgWoogIZ7oiuieLk8DYhURyqZvImVzO6NI/xwj1eY5sxivH2Lcce/XKORbjFPnqnvUzws3XbOem9vc//KhdPHrQ5o8etvX8Mcsqx+0m5MsehM7VknWQxDQ5h6a7uSzQ+bdasl9XROdJ/kBaYYtRlUtIF7RkXy3JsSl7ik3bvfNV+5Dr6mDCaZiQPmxWL9Ey2oNMpP+J5BoEzeGhUWSQb+IRYDjW1CHqKgln8sHYos24Eealnc5VMZbg8r1sz++pxh5TKJdwZpeuwM699uKdts4TMaS7Tf+pBjsMGjEmuYo+2lmRYjGOgTHl4GK/RmDV3nyhi1rTrzqqj3PDWaONS04tdVP+1DPziNgKsnB394zINLQjgm15AQ7Itt/JQHhJbDWWYvqxT8FvxLxfnDEu7jWmjcxpxzsJMex0bIychGTzWUUcy11OFc0At9Fo7aZoErzkz3anU/ZfOz48PDymqoDxn/qDEnPRFNOc+zC9NnfLnGM9dQQ6At8eAf8e9NQR6Ah0BDoCHYGOQEegI9AR+KQioN/nhWetnzfee/65F1/kJL6X8HEPdGzD8eUHcox9v1kWNzibeUpjuo3l5GukDrBtIogkvW6zS048+1NtrB/O9FDHMtvbV12VZ36lKENl80rW0/WqvvcgKrh7amLpmO2uZfiu02/yueSGHEkeriAsfB7qhO7pQwcRoV62k1zQefd9O21kSh3giFeqfN/tL5d+6r9ne6OWKpVdkg665mdsTh7OPnpZTxIt2g1Rddpusp3LH2O5nXo+oRukDO8hmygd17gWOSN61R7BghP1IlpLIoRku9j/S9xiqST9xLJBylDSCJ7oG/3ETHLPkxcP9mft6JBdsdA1lhkGlvRNm9I7Ohj6KGLUvJo3Ptv/9mWeKfoG5/PHZ+3xo5N2cv9eO3t0vx2gxwHLGXeYqCP0IO6OOcspiiLK5JecCzuQseJkyiR+odAoWxKd5Mo+W81Z8nfG9Xg9ax+dr9vllD25dvfZkH+XZZdEjjEPYt5AxhjhdOMGEWVx0mLilnMxl0Kqr/Og5kKMhZlDckzNs7zKqm60G8bZ6hI8jpsEquNISzM3beudwphD8c64r2nntPTdr70w9tkro8yqjHniNyG5Slks3xz6e1rHnKlpnxFfjqORdDdv3mw3jm/GSZX2tcNecGEb5eIVaSADLXd/NvN3ODzB/cR2wXmfZatOw+lAOEqUSYzZj8kpG8ucJQ0hzsARLcdjn6Pe5XKPMX3hD/z4T7zw+g/9MBviOTYxPvzkx+43BVSpW0jtPx2BjsB3i0B8Vd9to16/I9AR6Ah0BDoCHYGOQEegI/BbR2Dj3KUInDp9449JT5fuPjw5fZHoqBdZorSrYzmkMWQMPm0uTXJzezxN44bCATfyKBz0LefedpIKle/KPDcS971In02ZdfU+SRExxaORPEnSJPFhXdOm3mCTSxErL6ghyIDBuY36/kgVWCZpV3WNhnNzb8tGFOj4R+QY9e0r/oc8AKgHG3pH2QKnW0ffyKVKVzjZ1i+5eU/gMt/oKvpQ/cHRNx8UUIZ+LPMxNKFXy7hMRU5EJA8tjAAy6E2MkoBs7f79x+3B/RMrg1fQPBtdoh90Vt1YugdxJRIbfQYCjQYRlSTeYZrvw3hsSJVhLNUUNYJM2ybYqn7ojlw3T3epZNijDpI7RmKhuxhKYkh03Lp52PaJBLIde94xrSjVfupJRiXNk3hLZkjcSP4EWaLNQ7J/L0Yir80Qie9VO330qN376IN2/6MPiWJbsOfYTrt9eAQ5Biac4rgmCk9pa56dF6E7+qwhxyTvtMP7Yn7J3liXzAv20SIi6Xyy1+az43Y6PmqnbIW/nhEVhVz3rRNCbSxdDw73IARZXrm/SxnyAuM8nKD0N1ubtWMsUTkkMQn7KHcM6jtRduT7DXLFCaOWa//wTubm3WfgiDbZp1iiK33ZxrERZ8skk907TWLM/uNislpnO4VuEo1etAl9/Na5apmtNk3px7p+/xP3E4Mo3GMPsgNOMd092GcJpXuzgRnTZG8P243eYg6IYUTcUX9neBbLQ+aO0Xi7cXLlLAi3IIixUXIsIs80dogCs+/4liDI3KuN79oN+V2NyVEGs5dvP/Pca3/77/yvx3/4j/7R0JOfsCVsBcsQRV5PHYGOwG8Ngeu/2L+19r1VR6Aj0BHoCHQEOgIdgY5AR+B7jQD/m9X/2co1Gu+/+OKLL+FYvoTruK+jOyTcQzkCImt0vgcnMRzjwSEux9j6PtfeZNb3KllRtkVsWL/k+GyquubXVXk6116VH/W3HNmqt7kP/qz1PaXS/CKeqq+QNZAD5m2nqCsrFTYYRSOJkElZpcc1wZalVW9DBg7yrV+pnkuGdZUp1kFS4JFbVv0U0WL7ssH9x+YsWwxmgXzrV5/WM7/68TWe9fSHvoIIGjANhgSWJDZkjzlhC0UkUSMpt51qvy+JlSBskBtEIJXUGSuSXCrAqrE2Ws58OoIw2iHyB24uUuJt25KROj+Ng+ViZP3Cp+zcfte++Tn7gj08aeePTtv88XmbIX7Pzc9iWaM6QvYiZ4Lykr+epLlecvokWFa/8DSctriIfbIusXPpCaH7N9veMy+20Y1n23r/RpscHWf0GLLdn0v9HIsJ5JPLACPyCWJOssjvw6Su1oEXjL62x7j6LrtqXAM72tYcUE6MjUQeyXIvy7dtqL4qLyrzs/2eSwrz+yo5STrVd58Dta2Tz5JR1q/kc8n1ru1+OT5bpm5GixlJaBTYAQTZlGdJs13IRceGKrGs26/O+rZzj7Mdl6dyHbDskmWRcR0f3wg5yprFPmNE+EGSzefzwDfHAqKW/j1cIdMY3pZzeRnbxXJ9xGf0xnPPv/Dpn/0zf5aN1qgxmlA9QgBDxrZ9g4B+6wh0BL4LBPL/knwXDXrVjkBHoCPQEegIdAQ6Ah2BjsA/HgJPsRFPkRpPycajxfM0UkXndmd/bzbdfRGn8SUcwz0jp/AMdfRjn20qhYNZjrkLlYIcwZuMO86nchRVS9J0SE3s+hNt6Y9nKkTeQJTwXPXMr2fvVdd8k++RB0lhlI77HSGZOzpI43G5J1lE4tC1MmJ5InuBubdVnRoZp/gFFYVQCTBgQzIRcQUYciwaIsTcxF9ZpRtvqrPRR8IjczJKRhrBuuuBVRqxIX2KNjpNUsS2SInNxZAb74mLctV5Q4goeMBMLWNDf6ruQhCcQ/zo/IdACSmJBHUlLEacNlFeRALFO/0pKjDiwagf95yKMjumXkSYiaPtUVod1T300TB0M3SQktArxiPaIq+YruE9SBpl+U6qfgIbxu6YSKA9xHFEKtPQze/dg4ramsI/d/qKfphg/jPczrbuVaYsx967+79FEkjr2SH5YvPw/v12dnraLk5P4mTDHfpZLS5jD67ZDnu5sVSSDMivZdvbDwNTlBFjiiGkyY36L/0WIMZWvE8PbrTZM89Bjt1p89Wk7U3ZAH41bmcP2d8MvV2qa7STEYImo6eMWlTjIGrBMPQWY+Zl4Eupp2eqeiw3ZR47n8XQby3scp5j/xAGFmMUmJpHirJ4ymfLMj/lXPfJ3KRfO8sq4mib6+9TWXUpI8aS/j2oQIgjj4cYF3+RlVpYzDg47sxD04rlq6oY/QMxAWTsOTYGb6Lu1keQvBzHSv2PPsylkRJqkphXzAdRcx6LyYy/VZJkM+qKo3NSwuwSklVyzAixU8Z6Pl/E2F9eXgY5qQzxdxxsnzi4VHY5uuKUgckOy3zHk5c5AfNHX3vt019mMv4jOj23HktttVaNCaMVozCp/3QEOgLfJQL+de2pI9AR6Ah0BDoCHYGOQEegI/CJQ0DHj5SOnx4fO3b/6I/9+MHewf6rOKOvULZLHdmGNY4xj+EaBnFjw23H2UomHWhTlUUT3usehUN5PdfdNpWqfsmpu+XhpA91I/qJPIkm84uUs33J2CaaSk7JqHfv1abu5pnqnhEoZSmg4Jh/s3a2qb6rvfWsv1nCCerbdaxnKpk+W56kyLUO5ilL/eu69+BRuyCyCUqFK8mNqrPpI4buGl/LK20/w7ZAmDGGkA+bQxeGMY36OVuyKXUyL3WqZ+/KDEIjphfvEniQT+ZrI5am/jAqz966AbmE3pA1pYt1EovEu/IZ5s3807ayr3CzXsyDKqP5mn3a5ueX7cEHH7EB/Nwd2DkgIff8yrpikf1JyjhfXGLpvl1uqG8deWJpmqWRdG6+v3PYdo7vRARZ2ztqEy9Oq9zdZ6kg+2HVOJd+yjVSSlmzIGhyHzbLE4/8buxbG8yvu3h+s2Sdkh/4YJME1RN5Ww2tE/XIq2dtzOece0G0DuXKedoOxV23SXnWK3lpi7VSD/O3y7Mkv+HCJDbqhyQ7YpmlyyWP2KPtiKgwl6EGqeiYwKblqa45TozOZpzFtTb7d9ml5NcBJ4Tmsku/Caeee5IRFejJq0Sm2X5JhCD2OonH6mmkGdedy/ny9//QZz77+37qX/5XjkHKTyKMxo4cJAX21BHoCPyWEOgRZL8l2HqjjkBHoCPQEegIdAQ6Ah2B3y4EcCVDFNTEEyJ1CjNBw6wn7Y988Yvtz/3cX7qJ0/gS+c9EVEscPBfrCz2LUY+cfXtc+oRMHHLfdYp1go3Q8N8KL11HPeogqBxk+4pnH0g6qepQEUDW992AK31So5dMtvGqZJ3tPCOHPPEw/Vj0wEz4jJAl0WPEUURJIVcCwqTORmHh/tpR5EkOpNwsTy0syv7LzurfsBQR1eYQM+hFxyFHcgHpxpzEu3YaAWNAjQTNtQ32X2Mj6ZC6Z1SXUWRJLFEp8ZGwGTDXnof3HhLlRvvxThA6IUmyCTInoscG/CIaDKbHUxjVqzB1AWyc5mkH1A37fMQ+obFcA69GLkszQ3uVkK8+S3Z4QqHjwLZODj4mQUioFtFa0afNI8O2EmUZ2ffcM8dETfFMHNdifhH9q4N1KtV+Xeoc80zISOLgOORyxiQsLTd5NwLt8vG8PfroIadXnrJGkigvIpB27Y9II4m71cxxIaKJDd+NSptOWQKJ/m78XmPkwmLOtmzj2V5b7xy03eO7nFR5Cwr5gCioGe0lwIzo222HRJa5tM9lqo79lH3XjEpcT5EC4RZRjmrmOGBn6Iup9uX7FcoYM2e0U+Av3tpDHe0tVPzGnGFVJ8dpwIT610RWNGfyu/+We7pd8zzRnySZUXnRxu95mL+OIynqxHj4faLHdfMnyovcu3KODbY47ixgzHpgoazimar+0dFBzB/1z78Bo/b48WOi74jS43JfsmzHeNK5+6I5H6SrlJ9LVc0DW+QfQLItl7Tl27i4uAhyTAgl0pynqBFRiYymhPqYfyO+/avxeDki2OxosTP7Xefzy9/z1//6X//7/9bPjt79H/67vykI9hh/kuzjyVSA5N/B31z+ZO3+1hH4nYxAfS2/kzHotncEOgIdgY5AR6Aj0BHoCHxyEdDlxaNt7Wf+1M+2119//QWc2+d0RE04e2scWRxDKgxLr9zQWyewnGCJMt913ou4qfJBRtQNGSE1yQDft/Nss31tlz+d/7T8IA50XL1Ikm/bskuW7bbTttyS4b1S1d/uz7LK3663LavKS4fon65d/mWZTrr9uMSt+rVOEgQZBSUxtjLiZejP8m3dKgLngw8+9EQDhtGInyQhbBN9O26k0IdxIneDi+Wh82BvjLn4mG8j5JnKFvMj1d0XI6ogWIzQUZ9NuXL8D5JFks4N+2Oje8iSCfNHPcyfQQbd4hRDFxXWYQvqEbqntNRxy67cIyvJziJZnK228wqi077RwYjCs9Pz9vgey1DPF22XmXG0Q3QRettGPGvvLNtqg3uQzSDJvNy4fg3xMoIYu9rl2jtkn7FnuW638eGttpjstDlDtIwNxEZBkHkyY0WLaYJy3S9L2UEODd+RBFeQY1YiWW/bbvNifMRySNvlPtdV5UmWiW+SzZuxI0eyLi7kBTZD+6gjB861XS5ltiHfqFuyvNez/ZYOlbfR0eBT8JfA8qp8747bmLE38suIOqO9jP46OjhkPtxod+7cIQrsANwYJ0lt1LONyfF3jLeTMsXPOspU3uHhQTs+PiIyjYg0SDij0HKMExufgYSm8V0xFdYcZDkaQ469DMf3hdnu5AvFkrGVAAAgAElEQVR/4S/+uzeCu55MYb8mBFUO38B251vPhcFWVn/sCHQEthDoEWRbYPTHjkBHoCPQEegIdAQ6Ah2B7z8C0DHRabl2g7vtqy465JgO6LS9+eavvvDqpz/7CgzGTYkDHUdYDX7SudWhjGQUyuAoZh3zqTMQKkZ36NQaORKd4FBXW+uXu2+UjBVomWK36q3svxSlTbSjvFIRI+aXIx+loXPWwv0d5NKHMqwQOuLgywdkg2hvRckK7baOjm5EpdFu2+kNOUPeNUZJFtLYjpCHPciWpDPZZilRRNxK2poEY2gHgWBETPRrZXCVOHBfNSOMjDjLfhLjJKEGctJu0PODDz6Q6QmMI0pMu/D8Y781SYAhokelLIpoMdqF+ZSrXzRR/yAj0HIz1gNQ1DEiKU0TI9olexI2GxUV5J8WUuZ4rxYX9EZ7I4gCCi0mn1MgFeUeaHsso9uLTeslD0FInLhHUqZECPXITILER0OHSNYTG9+ChEMfbXGPKpfeGn10cXLOxvyP2ynLUHeupm1fUgbihhWdbNTvPOakQxkuiK6ZBwVQHuRN2IArJ5mHsovYd2w3SLHpM3fb9OhOOyf/Epl58qbzhRWXO0Y7ub87Y03Il5vQm9yzyxNg1TnIxFliVLYKZRFAHhRgsqzmm++b72WwW91i7Hg3xd554sO788D5a6plkoRKDfOv6jgew/NQ1zF23sWcc1aQvxZvx4AUUWzkb/dbepYtdE11MPUjUwbd8BcAPBgr54H6meNea8hW/OgSfXeoe+MgcJs8vgBzyoZ553dQ8r3H3xOnlfK4GC7Khzr8fdpl77IRGC+X4yDa5pxQ6pzwmwxsaOjptCyizT7oy2nqfmXgP15Mx58+P1v9wTde/6F32u7slxB/GnNswSZzmVh2jmkBYfwM2f3WEegIfCsE6gP6VnV6WUegI9AR6Ah0BDoCHYGOQEfg+43A4FrqweLKTnYOZrPd13D2uVaHKjNE1rg/D7621QayZnCWdV5N7lVledbRUU3iIgqpozMbEVNUDyc/CrJetTGrnO4khFJ25W3Xs651tu/WC7JEr3VI5nmZQifdcvXUIyeVjJL99HvV2ZZjnvWL8PPdZF71lTnXv+bn5uy650mOhR7qwmXylMhqX3m+l9wqC1lDpJbPY4ibt99+FwG5nE+iJZJlW1gMuSq66TP6GXAcPP1rHciPPtUPWUVIlm7OBa+IEBtsqH6vIEcktkaDnoUrCqUayJNwmUJGGW11kwifWJpJFFol+7m2/ZpMqjzrVR3lFz6Vp75Bhlyu28m9R63NIcXYY28KobUz2WsHezc4AZFIL5dbgt3yci7PEuNknkSR1JvLJ1djNn6fsNzy8DhOqhwdHLclUWjLEdFj8MdLtn8TRvG2X6PHXJ5pJFPmSfRkufqpb+gMBmVPjZV2VB2fvaxrXiXrelV+1du0VW8mQsmpdpmX+ZVX5JltYzwH/SzPPJ80LnWpPqpcHSpl2TXBWbZZvq2/zxK92jBFrnjNILRiHzEixsTuxs3DmBvWy+i7gbyEPJTENNlfXjWnnQcSb6U7m/czBlOIMqPRIrJvjxhCxsi+vWvXEgIZO1xmOXbeujz2bH7x/MXF5T/17N1n/sm/8HM/d2vtIEeiIa2H5yGv3zoCHYHvFIEeQfadItXrdQQ6Ah2BjkBHoCPQEegI/PYgkP4jXumT4p561WW35konEwdw7/69k5fWq/FLtNtdQ1a4LMo1RTi0xFRYNaOUDLXQwZTswkXF0czIDfNM9hMnGfLgsxFe4X/zDFUQzrLL2Ew6y0XqGJ1icvHUtkOdjveTBJR9WSd0N+oIR90T7bzbWZQNsl02RmHINqpqVE49+Vqw6YtqRkEZHRd52qU+5JnUvQiBupcO6hF4DIaGXmG3bdIwl6aaXCJm+7IryKShHWgA70CcDPZxi2T9SrWfkiTmfU5o1GcPnVnKOGYvLZMRM2XboAG5uTQN/kfD6M1/pMAn5RvA5JiEjcKG3iuj0KoPcAiMbTeMo++bhP5GCxmpk1NswA8iKjb+Z+mo+ir/zjPPRuTW1YoTJR0XOhaP0Fsl0IWqdhRzLrFDl8jKcZpAYtlW2UF8uJyRviTFzolEevjB/ba6gCxZS3xhLwcS7kCCHe2wP9l6DiKXcdqk82J3lhvDzyDAOLcVu4kQg0gbHdxsq73jNj643RajXSICx21BxJLzKfALUz2BEkInc+IbcJxcOqpezoPQk/KwFQov87M8xtf98vwHdvHNcadW4DHlOe3M+ptIL+sOk0R5tYw39QqkotzvMOvZHmhpI8SmmAViQ577qUXZIDPbiLlRVyE1xsi+Qg46i73zpuY0oxZTovpw3BjBmDcSVrar+azcMSTkmvkooWUbT7iU4HTjfD9f6xtZ5x5x/l2axN8jdXFu+Z0acZk4lQ5+biDNj3WugmgTPyMLF4aLmYvwMZ2RTzNPJBlz6Cb3q/HeYtneOD2Zf+Y//o/+6i1Oevj6f/af/Kc2ETFqXP8tMLOnjkBH4DtDgE+5p45AR6Aj0BHoCHQEOgIdgY7AJw4BHT22RNIZHrVXPv3ZvZ/8yT/0En7sSziL+zqSQ8LvHMMdJNkSDi/OaZXrKD6dog5Obt0t91kH1nYR2cN7pZJR96fz610ZpqfrmVd9lVTr6PzHHX0tT53TifbdsrJDGabK334u2U/XtX3IR1bJr7retdfk3Xqmuvtsne20/b4tt2RW//GOPPcbm0OIPbhPhJSyBiLOeuuB1Av56jH0H3eYyFySuNV/6JJ22EYyTMIjbLBsaF82RX9RMTEASFulHj5RP2y1He3dC2wjy3aQZJIcxzdutl0Ii9Ggr7qX7RJlZXM0oY22lw6FV93Nr0sZqnR6/7SdPTyPyLEx0WOjJcslL67i2hlx+iGE1h79G8m0v0e0EazKlGWSI0g3N+S/2mHD99lBu5wdQZLdZg+yG21O5Nj54qpdzBfRR5FM6qguRj1J9LhhfyyTHSKWUrecBzFG2iqZiK4SSGWH73Up0+ftpBzrelWZd99LrvWrTt0juiqmQrbd1tv61af1k3gy1+TY5vdf/UX21o/5wf9CMdm+6tU36LtS1d3Irag/PHOjDQcYxBLX3EMsCeBx7CVm5NcekWVGkomncNheeyLRZybnzvUcLrsty/oScWBH+yl9+SyBO5Qx5ePv05qIsuWCaDJOhn2Bgyc+zSf22r/zb/95+EnqxlehiU+OSckfFOm3jkBH4GMQ6BFkHwNMz+4IdAQ6Ah2BjkBHoCPQEfgeITD4jd9GOh4euxbhoP+xP/Gz7U/+6T+7d+P49guXi/ULEBO7RpsYFYLDTcDG6MqNtIusqM3Un3QRrx1yIzxwIXE8kxAbV7TYEHmmm2lKRxznVZIg3u2VZPPMCOc1spQ5pO1IsyAEbIWjG6Em1NFZNa4n9iQKAiIbXjvM6VCXW20wlWW2C+cdBXSWfQ+bKTNVBFXpbV443JRXe6OEdOJNtq1y5WZkVPaaspVL26jr8kIc9vjNvleD479a5dJDMZlE6BcEA7KNVjphfy1P/GMtoEaoeei5lqjwuEzThkCQieA97JFM8JUMZJZtRuiUzeoY0XfaE20kZpRHX9GYF1kol6pZNwotz3GPPcssl1xBrzUnpeYmVkYA0SekyA2WVwY2iyECiJMWlyyLjLHYwtFldSV+bRRcQCVOaa+EX0QWEQk3gfSdEgWlHWcnZ+x5ltFjYzAaQ8SNCA1ankHU3thhTzLIr9VjllvyTKTY7j4k2d5+u5rtECFGpBF7ky13brTx0TOxvHLNUstzluBdMs5io+lYxg8HFUDoRUIHIyiTzBm+AckY0aZ/I/ucr+qnnX4efhPih/a0G8QgvOo4jyRAYy+umF4ORKbCvfBRpinGj8zruXk9jyyvSMmQzXtGeVnic34Pzp0RS1OjD6MCoyx1Xa0X0YexXlE+EFaOSdYnf7Axpg3j7Ripl31u9ESm5sXS1qyI8hwJirzFgog4DkAYcxJoLMvkRNTUF12I4PNZvZ1jwq/MlOudtmZSbp4Rje57Rs+MVeLiWxDL2BsnfI7jrwsBtMt2ORnNFpeTN87nV7/rra98/Vf5W/kVm9KLAHkTaAQN34XzoKeOQEfgWyIw/Hn7lnV6YUegI9AR6Ah0BDoCHYGOQEfgB4AAXjqRMv/6n/yZ9uzdFw9wU1/CkXwRRXbY2N01R2xEnf9zNkgTCsLx3bqXA68DGnUGMqbqhWM6ONv1bFmVa3Q9l9NsPZ3Y7b51dKu9bUy+m7blmZfkWDr4vquXdUpetYnG/JSc7fJ6tszL99Kz2m3LKRnm2V/1GZhsN+BZQkh5XiVbMqn62q5u+40u+OTh8FNBZ9/ov9Oz87ZgY/Hqf6OjJAzwhHzIotwwfZCsc18JOaZYmjpEaEmWYWySlFXPOhJWEAyRlCEuMkQm5VTUmidWcl3FUkrK1IXxW3M5rqbYqB4Cw0geN7NXT4kj7fXZuzghdINT2Wh77Sxsa25scKJcmmN5sWofvXe/TVgmOWZJpNFjawiXS/LnpwuiyNjMnZMqb3By4uH+ERFKLK/cYakfuM4h8y4ZkzlL/2Lvsd2DtprutTks5QLCSILFvati+a2EmPaTnHvSSDW2mZ/EiYSZ+UZa5TjlnMLU3zS3bFdjrVzfxaP68V7PlldSrpdl2UfKrrztdtvPLlE0hUxJMcckuKLMi3zKC/Nqq1zzKj+E8FNjkWOY79ttSh/rM9pMKzFM3EpvSVFJsSmRY0bjSSQmrtffcpJ01zZX/95Lp9LdPJ/Nl8srfXy3z8EWl5SPPZX08nLZHj0+e+Hs/PJHn3/+5c+zUdqNnL7xDcD++aH01BHoCHw3CPSP5rtBq9ftCHQEOgIdgY5AR6Aj0BH4PiHA/0w1Egjn/Dd+48s4h6ubOPvPLVbLW5IXOIl6zASRBZkSm/S7rMj3IS8ceJ91UnWwq8y7zmfV06mt53BQ4RLcV8gr9zYbHNehnX65VyzLGxxZZZTDa7sgwSRihhTycexDl6f6t0+ThIP1cnkUDrnRXhv5kBd4v15V3zY+1+V72VFyCpNysr1DYwzLSK2PDH/I1zFQlm21R8LEzfvj9MbQS92wKbx36lA/Nvcf6odeRi5BJOWm/uP20Yf32hUEWekVuoZNjK19DYRNOPbCIBbaRNQLKKNgYsNLKBsRP/JSA+mzsV1yTHnYQeeQFbQN4ivJhXimX4Twn4wPl8/om4n22LaWNMMelzLKtR2wrNE+Cj9Nt03ceQxSqEg53q2bmF+Pi0SK+epl9JhRVquLZXv43r22OJm3A5ZK7rBvGAsqIcswjv3W2fKszc8WIDBrh7s3IMoohxwbc2exn9uXteXUjflvtsXuPvuQsdQS2aysDFKscIl+3YsM3WIug5NRYtoeZTyJs+Pje4y7xB82LSTYGBjLhFUMrudo1r+WQbkyByy28zfPyHP++C1uvkmeneRXEtcD8aWkWooYfXviJEk5nnhautf3Ue2sq/6+e21sYrBCLSO6JGPFwOkCDo531EOqe5vlvMu+7DOTp03mwQ6rlSceYGfMA78PyDGi+Zx+RpjF90mjDak2TC/ngNGP5tflu3qpszowQJC0ik8SU7zDDqUyttbhcjn5RKz9LlHl6PHp+eeOb93+XbP9gyOsuFZaNZBZ/VVBv3cEOgIfjwCfZE8dgY5AR6Aj0BHoCHQEOgIdgU8cAumCEqFxcvKYkypHz6+WV3d1GsNxxHPURVTrwXEMA3SiyyE3vzaw9zmiRXQYJSuGdt/sXuVRafix/XZdn7f7ikJ+ntal3qtuRaz4XmW29bnqlCzfw9knw+ckrVJ/34OcGfJtU+V1j/bkb/dTzrgYiuA1nkP7rb6C/Brk21dwD7wHFSLRIVlGUuYk8pMwMs8+3YPs3Q8+DKLKTc2L9KjyEcvRglmg7ibSS8IEYkuiSxkyALAyAyEVQmweyXKJgiA7VM403LW97De73pPYQKZ2OaRkRN+SEfQrWei7JJI677D/l/3YXmIr2g/yCjtxcJ5Zx7qFf/UbmNPZRgeI3+Xlqn31y19vM5eewmpdsWxz4vOSjeAnkGBEBy3MIypshA6QH7CRuxE5dgEJcg5xttw5hBg7auvZPvmjdgEhuxQ79PaqsYZUjmgyeBbN3qTSs+xLfVNPCauyZzvfvO1k2+0rv80c/+3nqEPTkllyzFcP07BkOp6r3Hs9b5ZOhw7beKZO23V9LrnVPvpwnEn2G3Wgj0zbdaqddbRBwtdxr/dowI/1jCDz26i7c7y+cetZR9nbl/nKKh18rzbOIwlWU+nhc2GJHAkyK5hF0ONq7/Ly8g00/PRP/qF/4SaWUOQVoKYg3nrqCHQEvjME+h5k3xlOvVZHoCPQEegIdAQ6Ah2BjsD3BwGdOqkLGZh2tViMHj549CJL/F7F+by1JBosIyeM8sH5hHhYQyqkw5mRJkZmmII4wTnN2CiF4ozznhE0RozoRrJpDyRMObK2i8iUqBde8ROOquXqZSpFfZaosdttR9g9g8ISytXvOtknpE9E82Q7y6pO2qJO9mFdTy9kY3Z0MtXdZx1rPeXKs63PufwtCRvrmSyLCCAESw75rt0RKYcMSS7bzszjXaIo5BrZhoUCGvtrpTj0h+hZ5kbwJR+FaKutkgc77dEjNuhHnn2ZarmiuIjzkI2nT2QOiRGNcRPMK8NpwubBDsgDG1SUT+iuWEhPl3TyEPral2SL0UzeK0V0WdQjB/uCKrGOFdBRbs45Mp1CcgTekhVJkoibp6F6uunKSJ9ob6ScBEj24BwIwg8rnFcL5qqTRJmOk3vdOZ7G712cXbaTDx62MZFii3OWdsayyEuWWmZUE4xwO79cNDZib7ODGUsnxWfMfdzOV7O2InJsdHgLguywXUGcLZG6cCxSFTUh8Tvo75sb8zvnphB0Nd+1r2ysvKEl+QBCwtRN/VzWmAbbrpJtt9/NrzlZdaIfmm7qSlZTWBF3YhZJuV7Dd3wtJ8t9r7zok7qRN0RP1X51kqvu8+XXGbaBn/Xd1zDaU2afV8y9kOx8j/F0zIc95ySsKJW4WhPJZuSbeJiMChNj50W9x/5m8ea8yHL18IOzmXkbnPjwlB2ThF/O4lXcUJ77k8WebkJBuzHLzWkrB+f8W19NJuur0WRnPJs9i00v/ZW/8lfvvvrKK+2/+c//GtLs1M/C/njqqSPQEfiOEMiv+Tuq2it1BDoCHYGOQEegI9AR6Ah0BL7nCOgx+r9Rw8HjfvDss3dfhzf41OVyccPeB0ceDgGXcvD+6v6EA2plkmRGEhc8Iz2c3cHLtZ1tTD7X+9Pyqsx6Vd/nkO3DU2k7v2Rut/PZOgMH8ERry+rSVi9TySndKi/IF+p496q23gesNu1ta79LySaSxI/vT8u0XeZLklgXXWXVuL/33jvtS196sz188GHb2+U0RYZKMiX6H7B0SZoyzk5OYRKQBcQSlhJZkoMm5UcSBG3Gp8+81CeWSVpBmZI1g2x1DiJCoeQVPlYNEiyaQAyUfPOxO+kYa5HQzQg2MaJTK+SsQ5fAhD4kUyXEbFtk24q66ljYKipxyrlTOLp0r8bBOtfPjCVc1/137rWL04u2nkPIQeygSfa3FZE0g9BaMZ5X7D12SVTZI0i0+8BwTuTYEnJsCTl2wdI7N+RfSKwNutifSV2G5cjDe41lvMbPtV6Z59LYmjOWKWOzRJQq5mlvjlP2UXnW9fK9ku+mKIOMUvZ2XpVFpaFePT99V+627Hrezq+xqby6K2vbrmpb+VXme5U5D7wWHHogjl5VvyLGPM3See+9ZNS9MMrvJuWW7crxeygszc/6EmubZZKMaeJZda2nTh7AQH0kuN8cR16Mxi/dufPcZ7/4xS8+z1Ti3xhlx/DDgf/1gIQF/acj0BH4OAR6BNnHIdPzOwIdgY5AR6Aj0BHoCHQEfhAI6PTho0qX6NeNDy6X89d5eB3Hc3/NCX86h/AYnFmXREstSTKyKJbx4YivgwBKBz+iSJCmqxjOK066yQWabr6Nx75x2iPfbrkkLXQwdZi929a7csyLKCXLeJd88QQ6ndyMiMH51b1FTrWPtsrDoaYSbXSEk2yRYBoTkWWd6BepRhzFRbUgvuhIWfy3kVmEmE6zZSYj5NQ1He5sm3s3JblRehgXFjbpcGtXyFaGNtiH0mjD3UiWJUTBL/7iL7Z79z9oX3nrN9rZo5P2hS98of3EP/PPtR1OVoxoF+obUSMmLlk8PYUgEzdkuP8T1g5y0ZN+lR8sIeTbBicJqAHrUIRWjoYNXQKpLPXNssQsxLAHVORDwMXddipiXU4ZjDx0gpGKvBH6RJ7TgTpjN+SXkKKOtgcRMUQ1oZKwkJdzReJCMYExbUN3bQy9rZwpxxW7MXXMmk22dG+nHzxqb/4/v8q+YzsIyEjIK+a1nV6xHHIFuTbbRSk2fx+xt9g5fc1pfwKztto7bHu377Tl3g3eppA2dGr8GHqLv3hqU4292Ev0OU+yjPriSN2q4zdDtbRBHLTDWcg4xpxyXgoIuZ7YGLLUFViDqGS+1dyjEvn5Ts/xHdY34MDZJk4eteKQ1DfwA9uQZ/8oJG8a4xN9UUZ764Xe6sNlNJ5Wm1ZhB30yfrYPQ8ivuVT98KGGHL9ZZUkKmrTQ+eLm9+avWbIadzKjLWVx4i3YqUfoSJ9GSlqP4qhXxGwMR0qN+mELH5N3a0fEHHJCNvX8++U8C4yiL+YnSvm3zKg39XQ+2TekW3yYknZ5gEZ77uxi9Xt/+Zd/+UuIOqPyiVuxoUvBo0QtJF3Pz3zvvx2BjkAh0AmyQqLfOwIdgY5AR6Aj0BHoCHQEPgkI6KfiAeLQ4wO+8PobBz/6o7/vNfZRenW5WO1LWgwJ/9QgMvw+HUau4EN0PsNBz1qWu3SwXMJ0RrPMNvFuW9L2s86vREmlqut79FUF3Kudd1PV1Wk2Vb7POvTmW8eArHCs5S4ima/bnvZYJ6+UEc459UI3+qry6p9alHrZLgRG3RWki20k4MSvMCw9cP83eZ7aaF1lmyRPdom0Or943P72z/98e/PNX203j2+0i4uzdnZ22v7W3/ofWdq3aj/5z/9hyMZd9syaqSCkGpFiOO/sj6SRQaokoaj8geRA1QmyXTIr+ZEkXuqdfTM+Pogr6owgB6447VEcQneJm6G6Oqfd13KSGBmAkCCVQIEoKmK17JfIU/7YPdFIsSwT/cViJklVYFIm1pIWORY5BtGIH+uJrfcYkwHzwBNywvEer0bt7bfebg/ee9AORvvx7rkAbCxFO+zCotGEOXu42/bAebXPyZSTZTtThxu3287tjBw7DzJYW0i0dbnxEnwkybSr9AjdSx9lkMqe63lznRcV+Ak8wQyBlZU2Id92kQa5jmfZbP7T8p1f5vlP3Spt9+9zkNUUBiHEe7Swj2rAvfqusVNPJVa+VQPvQTffTaGf9vg8kJ62sa73ah/fB38/VhCW9uHleNv+mmgsgsy+cs6EHoMcZcU6SMY87C4IGbPr5d2Qjch+on/JM/9F+1zWqfFl64K5FcugySSP2cxk0h50YwI9O5tOf+/rb7zxa89zvffWWyfKIqmgD9fAm9tTR6Aj8E0R6ATZN4WlZ3YEOgIdgY5AR6Aj0BHoCHz/EHgisgFvbz02YuJf+uk/3v7NP/3n9m/eeuZlnMmXcBz3iJbAfeRUROkOXL5wDlE0HFxcxnBIda2RQsV418HUETXpUcZlBVI5oz6XrFhJuEWOWWay3PrRF+9GYFV+3rOOBIzRY1Jd9m2KfnSQbTPIIbwjZQ5yrAPnZ3Hk45Ejgfps3j4ZSAheKNOWrFe6hN1pcDj0KWtw0CGFgCZ04Ilgqoq0wvm3Taikrp7UVw5/KB1Ey4cffth+4Rf+fnvjtdfbq6+81B6fnUFsjTl9cTfaf+nXf73d+/D99uLLnKYIgbXDyY9TT1iU/ApC02gc1hXuQGgxrhzCl/1iaJZj5bApvH48lgnZVlJH0F7jukR0miQUJw6KI7WuJG24HDftiZMU6YcmAOklyZV9pr1kOh8Y41jGKUlCVmHmXCniosY8+QVIHAgj91hbGbkTe0LZ/zXRYrsYCweR5Oj7bncjxvHyfN6+/I/ebHBe5FPKnFjOmc9zTqwEr/Fk1Q6P99vt1263gxdvtuXBus2nEGBHnJR4eCNmPruSQY0gXxsdT6kScDZCbzkCGzGg3CtTzn/ngCSPKW3N+Wy9IGFi/qhStrdezpsEku5CJqhlFBm6h4UWkAL7TZ8WZb7z2DLjpkbgNwaHeLc/UkVwDbUZ4iSRrwRtk7BxqC/+YR96ZBZyaZxLE5WS89oxzZRy8rupPO8SVsTfMQ8iEgu7xVFiPO5Df86RmBMxmZiC2OASy4hxFbuhH22KbxrJhb956yDGnI9cqkc/7K4fdseyTcpz3vh9OGO01Xvpnfj5lnZbJWJlR/xdZLgYj/Vk/+pq8qkf+wN/8If+3v/5f938D//yf9D+xn/9Xypqg0KMFU176gh0BD4egU6QfTw2vaQj0BHoCHQEOgIdgY5AR+AHhQCO5x/5F3+qvfz6G8enj+cv4+6/gOvqCW4LnESdvinOp+/hNAbDQSauZb7rGVItquLB2kDfVIc1NubmnmLI3EqWRxSXjm/J/k3l6XPa3vqVNvVDvcy1PGWqw+CrDuXeqv3Tssx3o3YjnjaOMQ2ermcvGxlBDGQd66mPSaJOekJyLEgD+rW8ZNneS+Ih20gwsMgOYmA+h9D59Tfbqy+/0m7e5JA8nPsXXnwZqeuIDtvb3Wn7e3ttn3vojLISNUbHTCc77fHFOQqm3aknz/TjclSjabINjcSilkaiC8qF7psfbRlD1FhP8lISx0LqSS5oqbK0yUoSlBREHfP9V0vtJGwwlPIkYmxv3ys2xJ8QseUSwgWRb+Mg+iS8coyjH9plHy63zLlWEUmqUzrUPTCWCGMUxP89zRcAACAASURBVPaj9z9qj+8/bPtjNsyHZGPfd9SFkGHB8Dk677Ih/9Frz7bjN54jWmyvzW5xEVF2RkW3kvdAiQXirpcpSrYICv9BjpmmEDi1zNHIslpemSTM9Zx1vE1FBgWekZN21HcSS5rRUTRrzmiL7VOmw5BzSLtN3i2LZ+pKJlvCaOV4bXB07LJN1B3aVz/beXEYA+WWeZnUI8YFGUbhZaKM+SHmztOqY1noR5F351HYwbMYrB2PId979VF3cfSyPy9Ja+/u52f7mG0Qtbm8295M5IbhzMkgvcQ7MqLvsinxHPQPQpGm6BBpmH/5klOX35GEKkTaakIwGd/rDI1fvlyuPsUsufv7f/wn2t/4ryDIxCmhr+b93hHoCHwLBDpB9i3A6UUdgY5AR6Aj0BHoCHQEOgLfDwTKsY2+iI0gSgxS5Z333zOy4w6ExguLxWocjjyeIQ57MioDGRbObPjCOKwRTZQOsI5tOro6rddLuPQYM+no5lP42ziuRti4eEmCQQc46g4Ej/K8dIqVK4GlD2uxeZWMDrFAxz+aWseKQ8TQtsNuGyN+dLw3ETLkTQfnW99YAqb6Vk6RHxgV+q6QG7bmiita0yioIW4+oZ9EicpEvYE0COc9iAT1W1FnFk679U3SGu6b9dobn2rn5+dtZ5dlf5BGpxfziKDZ3U0sFhILtDk4ONBtT0JiNm5f/frX2pu//mX20tpFDpuYQ6JJsxipJjmRYyN42DSQNREFhD2BV6qRUUzaM2As1lavOhHBg9Ij9yBDZ4AMozWj6hTJpf3KoceQLu5Zh3ywvcQ2T3t0aeWMSLvZQIg49+RblO+qOslGl5Y63ybDHlYKDHxdHuxY01fsQeZeZ5K0kGEPP/ioXdFHnODpCZbs6WU00vTYJZX77eXPvtJe+dxLPO+03Zssr2Rczs/YfWxBz/TlWKunVJgHCDiXYmmmRBH9iY26BpHjoHDJy8SKZdplIiPmhwgpTj2lXKBYLOFFWcvA0eWbRhxK8FiXOpCbkjx8PdG/EXQpp+Rruktst8YxviXbS13SFj3jJFd6rDGKcY15MMgr8ss+kZd9YC/zJQkpIwPVU3uyz9CPPCOxQFxjgmQOMnCYY+5RZj1lePns5XervBXl3h1WcZwxr9TNyDFJQy/32fOLj78T2kMZK5mxLfVQnzjgATn8Z8WQ6XhVWnH6biwrju+bKkORcKrPABnSB/spr9M1nYzWI9qOQDvYVSYlcLfd8ewl8l555vadA0I5zwhZxCijQv2bVD33e0egI/BxCHSC7OOQ6fkdgY5AR6Aj0BHoCHQEOgLfTwTCjcTxg8sKb1JS5hau6os4lbfJwUEfPM3wH8ngNcmmbKojaj0dY31h393zy6TD6yVhYa4Oby650hlOh1TxPocQG20l25Zz6913U9x5DocWmVXmu89pSta1z3gPQgKnl/aRN3iukhBF5GQ9O7AXjAknuUi41EUiI0rpf0WEkWchKk9yo/oNOwfPu4gUZUa+TnaINJJGEg0nG7Ir/Gl7RL5RYDdu3AiiICNuWtvf2Q2S4ktvfhny5qwdHh62G8e3ISqSRFKmuNy796CdPiaCDE9f3199i5hKxcEgMAFP7wNxkfYO2KqHyiGPClwZ5VNsgv2IQtwZdJexZQQgbQZ8om10mPVyjzEFQ5JoL33HOIpd6MPY0c9otAcuzpds5wb1RgHtzPbA5aqdnN4PUjD6rr6oG/MEIktyJeTa3nLsOHnwsE13OXnyZE6UGhFrkGOzmwft9svPtk//nh9uz77yTBsfEdmGl3Z/cdEuLuftkqZXdQCByxohY1xoLF4mx0nx2+NmXo5xVIH8Eet83pSBXemXJflrnjbY3ginenZ+0kuMR+EkQRQkYGFIjdTHUXG+Y3aQlspWgdRVYiq/Z3HO+Rpzb3iO2jyb53jl8sm0N087RQ7/HB+X55rKlvyOlcmyVW3w4AP6c382LVCz6kvbLDNZ5nPgRt9JhOU35X50QToOdtqX9Z9M6MkcLALQOnFwBUzWRjcB4XJaaZPLbLUvxof6NTbe02564b/UXzK3/ubl3xL7Xy6gpYmudOkyYp9lyeVn7t597nVOtfzSh29/FRpWiwMfpqESeuoIdAQ+DoFOkH0cMj2/I9AR6Ah0BDoCHYGOQEfg+4wA1I6nV+rDXV3tcJrcS0TevISrvrfC2TXhpLszv45eRC3hxYYjm068DmaqHI6pZIJtIhQDt1VHGic0/UUrJoEVlZ76cTNsCZF0lu03BXsPp5v6Eg6+S8iEPlUHh1gnXXdcDsN+tx1ko8MqRTQY9UJ/ZcY/2kJWRXSKTv0gP8gA+qilcW5sz5tK0BdRPbSPZW/k2Z9RTnjZ6Jn96bgnv5K4XBM4EmQSFeOIIrPttT3jiHL6u//732v3iOh768tfjqiyw5uH7cd+7Mfa5z//+fb8cy/S9pqIlKDbgUR7BHl2KfmAXJN7bRHyApFDXXVCf+3O5XBR5fpHUoE66qGJEZFF5JA6xt5hLiNEREXXJXlDufurueu9xKgshITGMCcUHvLQz3/5POTRV6LkGHBRZ0oU3GyWp19KUEggnj9etPnZsv0ay06/8fYHnOD5E+145wgVOQhhkDkJQgQ9JezoPwgYIsiW7DN2sbxod15+rs0fnNDLuN2682x7/tOvtGdfvduOn4dkHC0gxIgau7iIJayOaRyuABE1xabVch5wGeVke9Rk3MVYnZ0FWD5EvfEYKaKprGioHf8Z8RW2o7XzRRwlYwwm1G73vypbKCI5ToZH5VuNm7jaV7Rnbo2MkqM9QxPjKjFmP5SkHiu/Yb4VXp2dtaTW7yPHwjFzsBK7aMSPMrUydXa8tN2Ud6yIbzLJurTHuvmd1pJrqg92Ky/mC80lpko/y2NJs9OTcTNyzOi+nSDHct8xe0UTfrkGe8NG5ylJ2exORvt89n34/MJu6xhNaHsOHvGV97gFZqkbOiFP4tZx8W+Z+kjOOt/V0XqqQCQfhSMOQV0T3YlK6/X+5ah96t6DR59+dP/BOwgqgmwSkX4Mb6ifXfbfjkBH4CkEOkH2FCD9tSPQEegIdAQ6Ah2BjkBH4AeCAD6fTp9uejj8+6++8tqrOIBc671gdlItOYCsa3UcyHAmaVvPdbLc4LPibidhFPKVER5p1s88nFHaSyBJ7gRpw13n/+m0kaGY6oDnyo87FpQu2+1Lz8qrNr777FUy1UHHWN/5iiiabV2u66TtOvbR3n5BR5ffOuMt0qraVB/hcNOH7+nMp61Vr3Sy37t377af+qmfau9+/Wvt//i7f7edcaLlZz/7mfZP/Ojvi+gyyQbJiTGb1rvcEDVC33vstbXkNED4zYEckBhI8kESpnTxbpI4ibGRefHRsZVAeyqFjtonccM9WyO3xmvAsSLDIjINraoegkO2YiWVkohg9MF5hQzl7+9OghBLHdXBa9L2WGZquadzfumtt9oPf+5z7fgYgkws/TfYomyT+eIrwfTo9HF75oW7bfYM8mevt6Ojo3Z895k2OULmPhv4Tzn1k2WbkmMryT0ImtxXi+gno/vYfCzlO2bMjQEa83wPXBhz77GEU2bG50GnIL60F72i7oBI1KeO/0zKSqIqXsOGyOcn7cm925TLyD/Rh/ViqXCU+UbK4cxnX9FJsnczHpBibtQvkehciihK6pRegS3yyOISg4qeGuYJ82WxYIc28iMNNwnuSMN8ihEKOYmJ2X7zprAFhYA55q5kaEaN+Xcg/xZYR538C2Vy7lUy38ukvhrnX5Qal2rrXUCqrn+K8lmlUy9xqHaWSeKtIU2DjOTd8tCX7qgHZzaOvRhd9jq/vNw/PDj41Je+9NanqPNLCH1gXZplB2T01BHoCHw8Ap0g+3hseklHoCPQEegIdAQ6Ah2BjsD3AoHyjK/9S3sxKowSQmMkdq7Ge9Ppzss49Z5eua/TGc7immMSST7HA86fy9d8V1w4loP8cvh1PMPhr34hDqIuLqzOYzi0oYDVkoTQtfZ0QB3YdDAHx518k/1tHHIcfOsYmuFdLmUN0YEALvuWzHAPNHtFHhEpUS/eSlY632aFLcgPA2nrUi/zqsx7kQbSHVpueSwJs0+9c3/zNugKiaJR5kcd+uHd6B0d68i3S8kR7UZeXeYdHB22H/78F9rnfs8XYnma1YjwC2ddHdRHB97rElvni8vm6ZehBJUnkGfuuYQWqbs60EfiQF/B9iT2vGU+cngk+aNeAw5iwRXjZjQOrKA2xWmWEQmXstU/5Md8UirEgxFmlwMQlEueuXfZmDFZXzJm8c5YEu1k28SVaCKJMcbUfbpmRJb90//sj7M/2Lo9C8Flvegn1OInDiBAtnoOySjGQ/YUm0whyIgx2t/fjaWpzo8V1xUblC0uFpBgECExfo4raEH6CMMSfEYGCxlFRrSayxrrlEfneeg5dBf9DuSoWU6DzEtC0XliZg67pdcpbBGXyMq54JiZghCSgJO/lkliokvWmJRv5JxpAp4ST4Gf82IoH43Yg453+4/5K5sL3p7yWGNpz7Yz+sx9viTSQlZggSTnptoNaoddyA+9ycv3xKP2EgvdJE9jPLmFXPRw3JTL/PQvT5xOCRkW5BiquQ+d89n5rWkxV4Y2ko1hJ/Y4FvZPjejfsWa0wm7tmrCPX+m5uUvmMbAVDZdLv/O7RlCkTV1lgLffq4aH/fHIM6qpvXuRyTkyl/YYk5f2d2cvzc9OiCmrpJEI6qkj0BH4lgh0guxbwtMLOwIdgY5AR6Aj0BHoCHQEvk8I6GHiNfIfDvPrP/KF/U9/5rMv4WC+DIETBFk40XqIeqL+DAREZPCsoxvONc/psFqLBum3R/10pOlDN1PmgRQOMm2Ul+VKzFRyEE1ZRq5Uv9v1ffZkRnX0WcfaTch95r9Bn9RxW7byrWPy7rsyol+JAwkBSIRw1FHCMsm2ahdNUTeizXhRhvZsp5C1lWF5ysFfRv52eUR2heN+3Ufps5A8ijIIG4iRyld795OaDXLFaQQhduL+YzIPOPeSHAIReufwpd0Wi4EEQ1ShDgRDYBLGDYr7PLwXaWRJynOzfA4Y2NTXfmyTCCIVrqriRuxGGKp7JfNcUus/50RGM11GHXFXitzCGUtGPYhgNGG5IySZ5NBkZ7bBT10CV/I9xdNTQCvPJah7B3txSTiZfzm+ZKornQWaRDu5fxq0H52hiXjwViaJeyQITe3PZPn1/Mk2zAXtoGERRBFZF/LoKbrLyCZl2Mar5k1iNYjnVvmZk/NGfeMgCnQxOZ+CKGMuiZdzyKRcy0ovv0PxcRycr9okkSQ2ceAF5JQtYz895NB5yFGGekhwmq736dOYTJs+tIUs60+R4V2Z2d66zC8Q8t3IQVPoSHe+RtQYMmYQpqm70yjrFU62re8tBDCeQZJBdLrMNKLjkCHxaqrvxGfnlpGKQfwNY6q8b5XsVxmOozirTtlr2zlRmjs8kMfbeEY03Z3Pff533331Mz9y8LVf/0dhMahGF2XDt+qvl3UEficjkF/772QEuu0dgY5AR6Aj0BHoCHQEOgLfXwTCg8XJo9drF9dH3fdR+6l/9Y+3v/Zf/Lf7x8e3XyAS63nIhl2pJlxDgyRGXtZMNzxV15k1lbPpMi+f67IsN8VOZ9N+ttvoOJbzWPciKiRwgsRBXtVLedmmnqtviZkghCgwbw2REBfMwHV+al9tlKs+vpde1pZUiPeI9NJyI1x08bnjKVtmnn3Wc8n0vv0cmFE1yAx0m0ACuMeSpIbRM0YzCeMleyMtQNoVait0XkDcXPKyxKH3OUigYB0gRogKc0+lIJLUDXmhD/JPTnKfLYmI0ION7WNfKrqiVQ6++OD0M7TCuEnKCDmUx0gLhAkdrojuMroPPhK5YIJ85Y4gZmiV9cTE6sPrlX1wyufIaD6flQvpkHcixli+GAQMedq3S8RY6IBk0wXLHh8+Om1f+erXUWHSHp6ct/v3HlLHgw2YnXSUywOHTd3F1DlGNzkGyDf0CnmG+qzWlyEfqgbCxMsTFY1ak8DRNn6ph7GhjzJG2iouCgUvbwQnxTywrySO7KfmqbrkkldtiLbih4y6nkTdWtspiTQJLfG1Q8x15CLFXlrYbbSkJK4kX155kMK1Hjk3nWNxOigDF8sWUV6iccwV0VvwSTPmyA6RWwaoORejHnfH2/fARz24ag6Yt6lLHzGVQ0tsdU7YPjPRnxcwmHEPWeLNZbaEpt+Qc9l5E98duDozxEDiz2dTkF4SgeIZczTxdVzq2yz7lePl97qdYn6TsVSu8pFd/drWPrxHj4xZkGPOa5Sxa+/Ijf0YLy4XVxDYa5fhXs6XN1597VPH/9Pf+d/2/8Sf+fPXA2aTQddtPfpzR6AjcI3Ak1/pdX5/6gh0BDoCHYGOQEegI9AR6Aj8ABAYty/+az/dXn3tjZuQMy/ivj6nI4lzuORe/jxeYqZv5/AFKUD7dEazeeWF87nlMPpumSfcmao8fNLwSJ90MK/LN+o80c5yU/Ydjwh48n9+ly6WWl9H2ry6Vx8ly3ohD6e+UsnYrmPZtgzfS1ZsTD7oZl4SXhAJ2o6dOuJGQHm3zEikvCRxJJCUBXEQcG5Fow19cKZeu2BD+vc//MhuceYH3LWNKzPzhpLxoDlbJoWuQ428oVuUD7LUW/02xBrlZb/3iEqC6CAzcLCfIuo2e5Vt9e1SPyOaRpA2niwpFi4ZlPiJfhg35X7prS+H3Y9Pz+PdvDoRMcfhyTEsGxJjl6S6UT0RaDBAdm97SSCT5GKOmWNyfbqj9a1nWY2pJI7PJvu1TpT7DNsj2VKXpIuXyYg1RG10Ny/1Tvx8rj5SrjWqj+tn9VFQzR3v5sXc2cyba3IvW+av8pOUzSWMRm3tcLJnbIjPXbMkgT0goTApe8tmJYW9VN7W2Xzfs76YJvkmCWZSx3ouPaYDqSZpZmSY5Jz9mkq2z4WhJJn5gQG4VxID87cv52fVrXz7refUp2SlpJhvJZQ7KKNI9mm2bQrvBcucF+DNwRfwvvyRDGL7ajpfrG5fzJeHn/2Rz4Uk++upI9AR+PYI9CWW3x6jXqMj0BHoCHQEOgIdgY5AR+B7gEC6rBvBvBoTs2aT8pM2X57fhpq4s1ivx3NOP5SPYeleMAIzPFh8xKAAJDsiOmhwRGEHwvmcbhxYSA482/APJQfoTl/ZKxxeC5TFlTwFzufgTBp1ojMqGUSLeNbRdNmjywDHkb/RP8p1XCXBbKHrbPzH03t/ZQsJpiQ1fLcfHWfvlYIAUDesLoc67sB0ZTTUUNfTLLWnHO+SZ9SaiuSySPTXgXc5GBUi8ivIknS21VRSQZHjEXtIUVfzlDlVOMnIMvVbRL9gwF1CwXYmI6lowUmS7DVF/gkRVwG8kVNiOuZESPKNuokEGeey1IhmIs8IHsmBxED0wnBVE6Bosu3oh11G8Ig5cmsJbNVx2afzoVKKMI8U447Mumdu9C21FMtEKY7xpOzRo0cRVXawt0/ZiBMD99rzzz/PaZ2QaUZ+GdVEPftwFg8zLeqyZRh3xhdbncGxBxzvyhY778pxL7iwX0GMjTjFeNPfGKFLhItN/OPuvlSpn7K1U8xMtKU9NJEdQ54oUHF0Th1lOnd9U2HUjbx4sIZwuuxRZa2vvMKRttCkUd92OVaSpOqa/Rs751yRaFK/mEMQTiIEXxV9Gv2FFLBgfzd7sR7RYy5/3f3/2Xt3ntuSbE1r3b7LvmXurMqqU1VHRZ9ulRpB6+DhgAEGaq+NRoKDCzYSBlJbGEg4/AgcXH5DtxoXYbQwQYCFBH1O1anMnXvv77YuPM87Yqw191e7WjiZiVQR315rzogYMW4Rc1WNN0fERMb+xFqDXenQ66Ls2LsVFb35fWAkusIz/mccd2krfUaG4zDMZRz/AYI6B/pB/3tGmICcdfWTLhl5cNJGdfO3Qg+XtyqbzOw01Bg+YLz30KiLz97VeC7MZo3PIQgI61UbnS/WxM41rD2lep53oEWfpNKXDEP94PmIXh1r8cUE6l9bhtUGRpxvZxbZ9YubL3Ycc/d4/xBavujT+Zaap7qf39MD0wNLD0yAbOmNeT89MD0wPTA9MD0wPTA9MD3wY3nA2DIR78PDwxvuf0HE/NZMJgNHA3aDSINDt6oJJBjYJiaEuIPGVr5pDW7drmap2FweHShWcEtoW7yhCZ8hJ4NGW/OzPxATNFCHpGVXrQLq0AsaQOF9BfohT8DtnW32dZFPyzE4tt9AXeSu+6TtbWMCEaFvFpA2P699b8aL/OTBP7YYjmAc/fSPYIpqeDZSl/CVlv4C2EqIOul7AQhBhTqzDELKZlcyrzgI/+HjQ87sisChX/Qp0hITfUq2dJ7LFJShev/gO+PVhx5B0c32usAxwJj15jr07WdtjW2CnOgKNBWdJUo71wanMrD9ha5PgAovdtfJPsLc0L1+83L1yCH6jvkX/+J/4aUFb1Y//for9HjKWVdmCglBKLdL+bAyoeSTQ+EDjlAZdNGFsYJJp5Gl1iBh7IXZkmfzjn1mvcGn5biu9eFmZD/pKV3v+V6W8IkMV4Tyqr2vPgfS9CeDXDkXkzLG7Cr1Vs/LeijQxbF5NgWHhm7SKCNZc2xPLVuLaXSnX7+2HtlWCWzmtl7bW45LNfRu1aVSW1ov9quvstTB/vh2hxcAk5fnorUc6QWznLg1oLDgmPLO9i/8Fh9Qr7HtkHqebKvts/CDnRxbh6xH14a+4Iesedu+YxyPYuT7HVprCzneK01bHGvx2mtEINLfAfU2k1Ee/mo87p9ev7y++hnXVyCkH+TA0EgLk/k1PTA98FkPTIDss26ZjdMD0wPTA9MD0wPTA9MD0wM/kAcM+wzchG24XO2e9ps/2x+2AmQvTycPS1eTA3FhBZiG9wlkzaioaJQgEnBAsi5my9CXw8ATWFZw20GmgWfOFRv0CToBUohOK5PMABueBpwe/h567i2IHXUD6wHE2M4IRRl0mzSVAH0ADI7vIo315tl9bufLeWcD0Iva3O+QGxoavDbAV1kmCi5ewkDKDLhGZor3dRYbugzvmG0VHoInqgT/WAXvg/bLTv0iixuKPMxS4bCp1Hc7g3FkxuGcUUbmmOeZKY+z+dmmuCUL8OPq7o7sFZlBF0xSnsPHYQSDzLn2MrbasC9+XtCqqOCZOsAsZ3NRd2z0wpbakgjIol3QIYrJx2/olkP/qWaLpXKGnYKvvR4iW4AQ3Xe0P7z/uHr68lVsUp3Xr1+uNq+3q9/97qvVP/1n/+Pq7/3d36z+nX/v3wVEEwhCD+w0ay7ZQ+ibN05il4BJAULOm+u3ssgEOekJf8/1ski7/Dg3fV6ac6Ybsh55UuTlG0i5weIqtl2RvXeSCUX8OIVnIbKpVA8ugEaxtltqXdXzFd4KG8VbnzdpUgagR2uAGs/1MpswU+ices/fnt2kgmmeM5Ysv0ofy3qLHQzw6hbBPM8w92oGpzyuPT9NmdpJ4fBBv/1CVl/tK70dKz+L4wSR3HL4JO4Omc9x5I7+NUCbY7K1kmuyx4bskhtW4aVLA0ynyQr/WEfSmdnVJf6krfzR7c45OqqbW2f90Rprb8PYei+vNpy5ZF58Hv0ToFZPi35srjyCsNHXrFt+OHY8hHW2HM/s/vTyw+HhL169/PIvUPJ/h4sPoyxaSio2zDI9MD1w8cAEyC6+mHfTA9MD0wPTA9MD0wPTA9MDP7wHDNj8dNx3+/XXv/jl48Phl8SCL8wcAyYwEBVbSHBnUGpYSEgZbTvIr8CepgEIpNMQkyDUALO3JLagBMEQdYaK4xNgE1R7fwlYUZBK0y+BtQBSIyg3ND9vgyP8LDp1HIAGeltskZ/F8X2fBr6UU/LV4Q9t1FWtS8YQfHewrp3yNJBOlkn0Lp4lS9lmgUED642+Qn/7pO9AvHWx3VJX6WoLZCZjADH2t77SiRd89+F9+MGczgL4AnA4JjY5f/pj+FUyFRq0+mzLWwAPglbS62P95xB0F905kT0T9Glt5ozbNyUtfpJZNmSzCZIJqq0BXAKSYWdK9KhbDEvmlfqrogfPc+I5DD14fp9tgPvj0+o3v/nN6tXLL1av3rwOkFrrpVcUOiXdsaVrjveuqxaJksqwVV35ZF0KoCz1GWqFxvXDeJ+EsYQyH02vhHpj5lhn0KtXzVH5o9a+UtUV38rQOxhqc+YdRr32zm2hr/UResCm3tqpDOmjU+ysuZeuzvED/GIb4BP+66yzo4CZGW6utTFe/2Tt6Y9ihu7wQh9t9C2StgsyKVPd4nfkeG+RTl/TDbcC85SzVfaGjFN4ZU6xvcdfsb7MgixfeW35YXn+Kp3keynle32o99UVP4z5Q5MQ9vxYsV+5sUf/q6dDUdi52Q87MnDQex974e/ZgDX/zDH0wsMCaC0D/iQKCgqiC78BD0+Pb26ud3/5/u7j/0oG2b/kBRYPeAeOR5E2JY+HgLtZpgemB84emADZ2RXzZnpgemB6YHpgemB6YHpgeuCH9IDBHUHdGWYxrCSIu/3w8f4XvJHtF2AaN8aNBpYGgCISYmQGjYZ6DjQgNoY34vNTAaPZPFTosNsxBRBQCYpiX5UErATGliGnMsioF68BOhB8Xopc6edi8K78yjKTB/QJ0M0UGZkz0BrQOsog9sSbFMMbA6yXHDoN0OXLxxJa6QlppbFeySdSYJN+GXRaqQfMxpHOshdIGiWU6Fby5Kee8ITmieA77fjX/BQBLutSWLwXQPGMrJPK5G2KpVP6ywXx3xVAlaDVu2+/yzgEyYE2iIIKUGVi6QTHpM9+0+1S11+SFgiSbWvqaSbREkDwoPsjh7kfrwJ6kL6GBHzjOBkIqsoX2+JRfYf+5RXkqwe+QOECqBjHIeeoJV/ACmS+ecmWTf0lUAadLx3YyQPdf/6Lr7OMXGPqyCWy5WdJlhxXfaxM+6GITuXX2m6oiq5kl6TtZupZUqfNxCmBrD2Tnte22n8UQgAAIABJREFUprtAlvOakbOQh5JgaDaX2Wzyk7/F9a/JkiTDiKt8L3oy7+h+Ac0ESuGF/nnIBKvCSREFZuEcZKCL02qna5T5POxpUDZnYTWtU2KG3yMHyruOPHx/C3DplktluFXauYNDMuYcZ71tlJeeBAJK27lde/n4MgWL7vP26Htu0UU/XAvG8fHcNFO13JJInl3ob6+vI995VLw+0FeRJUvXCMX54DtV/apu2q68zCcEAeAYb7anOqXdKyPZkOrw/FZ47ljpT4MTHB7OB7RWYao85ylrOUIEBMnazPqqeZNvnRPnmDzzAmRqenrck217On55vVv/W/cPD/8bTf8TPb+NMrVanJEJkOGsWaYHnntgAmTPPTLr0wPTA9MD0wPTA9MD0wPTAz+IBwwGKQZ1fogxDZJXt7/+9a//nC1Cf07DiwSM0BFUgnEZuppJYZBI0GggyVD/uhjKJ0zsBq6OK7Cq7mGW3iF/QfnpbZ8rZPQfHotxqSO3ePTVoFWwoQJ5A25LgCCu9kmfQNyIvOwKTY0reu+7SM+/M03O/Bpye0zpQMgLlfdm4zSPyKvImE75lg5mF+XMr2KdcT1GGu/9U1f1F+CzFE3zKTAuLy3QNj5PxN2erfQ3f/v7jM0kiaLU3IZHgKyRxdW6o1zmVM7xu3YPecpMdo57EfXpDoDDTBkBwLwBoYCa8IIWJcsexrcvWm9pPNCefLl2WGihjL0n+DEaMOcRsOdxdXt9E2BwDUChON4TGIDEwW7ltJgpaGlbgiulbUzcok86u1ynu/hFb1MPi6IXpBGxqTeGFqASHzgX6O8I687N2Te0JmMx/VQo9gl6BRyjHtvjw1qf6tk69zNTa774B8AJp/qKrPB3pRV/x9tutpZZY2CV+K3oe/3b7zxYvJLdFPpkeAmYkdSkLtaxqq40+IhYGiyTj8Vr39vHSi47BLQg0a9mXF1oacfBruMbzhrrzDp+RWS2uoJH/MB9QEOv2LXRVxSeqMxFy3SNm3mpLDiMr9JLqVnt8rRvFMfKM1lgrLErqB6VQb++jx+9H/Ttu2533am3dWmKX/kzz5N7TlmP9LNzGGjteLi6e7j/zfWLF39//fL129PHdwxiZFIc1XyW6YHpgc95YPzsfK5rtk0PTA9MD0wPTA9MD0wPTA9MD3zvHjBYAxMwGOXg6pdvbrn51eH49KvtZncrXEEh6nva8FUVgAGDYCJCegip+ZhNkdDUwJWA2cyUbM8kME1Wh7Gh7c/+368BZyJdRxPUGnga5AaQUS34eqh9olgp6TfQ9A2Xg7ACT7Ovoh2kBrHhW/RmfT0/6B5W52IwLH2CfXSwRM7imjYAgPCSnyoxJnSMMftIYK75LAPs5t9XaRqwKDn6T7kaIEhAPSlBgJCFEQx71JOMKsa3nB6vz8xwEeRwHv72d9/Ak8HiItB3UW+4BLAU7NIv1a/MCx2De0hkhUZai0iVPMw8o83sQDO9znLM6mK8HzNvoMindL3Iz5sfpYtTz5MXeScynjyT6qufvA3wY74NZ8anaHuSdbQtYgWAkDJkCgoKeshR0OrcTr11cK7l0yWrucfbiF0B8eQlXdY4HKl3OfOiIbPHeIv3vkHRrCSbpBMoq6VVz0a8MOT7rAjn5AqRulV2E1eeJ+XLo68bMvqUstTfteXbT6V3vJliXmuch/mrGfmJY60/3D+uPn64W73/7sPqm2/erd5/vFu9e/9h9Z627zj/zattD0/71f3jE4fOC1K5btFFffJhnl0D6OJa23L+mlf1yu+DxisVmXXV3/5q1Edfqp/AnmMkE4CW3o/nlwWQljeH67Xd1MLPr7NP0qKRwnXyKR1tca1I15/WTdl+ag1DA223ZQ7yW5aZSmag+jZN85TONVbZf5kTjnCr09o+4MOvvvrFz/67//5/ePNv//v/EEWQl1WJoFmmB6YHPusBf91mmR6YHpgemB6YHpgemB6YHpge+EE9YCBowEghQjTqN5Tcrf6Nv/zLFzcvX/yKcPWXZPFsAXL20LJj6ES8TxEkuYwNjwpcK1i1L0xDk9vzF6Nzr9wEoNRsG3qcrxKlbdBfaKvdPseFH1ezq2xrPi1HPgbaTdvtZzoJKJ9rb5lFUXIFwEKPy+ThFizHNmBFE8W+AgTOchZ2LNtqmxi2dIoRo+3vTBVqMqStdFQn7WkeXnOPWwW+NvBha2yQJMEOYZcgIwJlMqEvwBHNkbMI1h1vVXskra+eGxtcH9olURiEB8gYgN5VOAnerU+EN9oD6GVSjfyKp/XyC0zSpt8slY3IGFibQXQCCdux7e/FzW718pbtfchwiR4Aayxbt8ZR9Ef8f+Zb/FrexZ5aL45RB7cveg1QA4/2J7ckxAHYDL2KNzxxmi9k6GJ7l7ov/vLJumFI6+C1fIu8ISuZdzDIfGaOa3zpxly5pRJeigl/bqpecqVr/urRfaotMGa/JWNzt/xyE28VxwnUCiwLhPV5YG691Efq97B9YDqZX3TY0SYAa7vbKr3a3sCeXOV50aH10McX0NQ1mLkZ9PJxXAHMxQPmsrOSPvv9mDlW9/Thp/aDgLp/NeQy39IWTel56dcGJ1w/ScOzhS+KFr2jI9csKdeLN9AJkrFFu4tA2ZYXRchDWdKQPcaSZus0z9vNi5cv/+xXv775+//6P1j9z//8nzKeXysR6lmmB6YHPuuBCZB91i2zcXpgemB6YHpgemB6YHpgeuD79EAFcwsJhGx/9Z/+Z6v//L/4J6/uHk5fEzDffrzj/XNEtrwFj6O+rgTICPY7vGYsAWEO+uY2QTlB5SUgFZ4ZgSp0CYoXYWEH+aXBooOGyEGWg4w5zTCqwLXovHd8tmCFoAJjo1q3LTbv1qXHCgRYzu1DrME1BwilL2AGQbA8zAC6hMKOq3YPME8ADUO34cm/zp1SXzJqGC9IUPrQDy9pqhTYUTo0wHBp8wD2fWdDjUwZ34YovX8BE+RHwN5Qh352VgzizdZ7R+bPX//ut0NeXczW6qmT17Joc+lT1/Shr0BOtsaauiWYQJvzL6C14mB+8qSqTWcgW0wjb3Z05iOj7ApCpPkD9CgeEapAO+ADC7cBUpXU+1/9/OerL1+/Wh0+/BbgSgsFx5wDxyi6QIn2bdsl8OWf68fMs8Lzag31WhgMcumvrFHWmmed7dUls28eWa8/dEC2KjefrENfPsCfmUkQpE8dtwCFAZHwmVeL/vEtkSnobyaWFis7h+EjzWcqNgYoc40UedY1ayIzjz9qzmpNRg6ErlFFtU+8Oq70dNsoIJB/8tYc+vqZPh1qPR9Wj6UeY+W72d5lPbeMbM3EVnl3plr3eQUZWsivNRva+EfdLiCXNvj81ZyW3XEJVrZ9TqLjU+f56vbLeh7LyMWTIn/aRvolQ6uVenxBTR7q6jzL++Bz63oaPAJiSqNupRAz2/xr/AFf9xr0+T/yTMh3dw2ICGh2//gQkOzdu2/W9/f30cH+WaYHpgf+uAcmQPbHfTN7pgemB6YHpgemB6YHpgemB75HD4yg04gtUdt/9J/81ernv/rlF//n//F/va234AlKcDx5lQSXHul/DQAkIuN4g0cDUO+9GlDKLiNz/6kBFSBKU0FmB6rVXsFj+BK4C4B5P9TLvXR+bK8xdHPf8ou+eCuji+2la8m2vfkEJKA/GSV0F68CB5outAmIL3J7vDSOMfY16O4zwQTPrPup/rJP+i7yaD4Zq92DXr26r6+tq34W7JDWoF7gCCEBhNw+98SB7AMZclLCh4ZgVZih8VGh9faqn0uOYA7Agbz1da4hH1/MLsMDImwBLDz0yjWR7B6v8q4tfgUqdBvN2KSeMqhz6apeB84jz+12/D3e361+/rOvAPyg48+ijm2/ei19oh8stnVmn/X2e/wUvaQxi6zWlvT2ybdpCuQTjIMn/wLojbHytLQe3rceuQoODpDMuva6Uy9yTOSLuWWPPDK+qrn3y/biSUVADbCt5ofxwnXwbbu8nu/PHGoddlVAS56tM5BYeBwAPjWx5fmWScs5sxHerrETgJe+aVm7LS9QoAjkdbsZZ26DhFuu+nDreWMmxMHHN1aSijp4XOyRj/LqWvJdM64tZiZ9jtdyfnrOBc1ig31SekXD9GuPpe3NSzlYR+030UhlapvF9mXp8Ypt34QOOZlMrxTnYsvkSpPlT1t0Zb4E490q7RbRO7aodrH/ubzum9fpgekB89hnmR6YHpgemB6YHpgemB6YHpge+PE8YLRHhLfiLKLfbZ72918+PN3fHsgOEkS42uzWvpnRmNNtZuZFGU8KlHlYf4WkMMiNgakBoN8GkCNQp8GgsMABgmruE0gSVEvbAeMyeEzgfeY+aILsGGTDmGJwX2Mr6KxD75Va7R0gE0qnzQO6vVVm9DNQ5m5D8FxjKrBeE9hHXwVFGAEvDvDso7TDQMreqld2ARCgT5QyEwUaM4hi57DDtqqXftYtOSuMq6BCziIrZ4bWOWg7nIP0ZyYYAH/PHZOnf4Jk0t8/cYYUWWQpZjfFhqIvmeghuEGTvC3SRB2MUavoNLbFUfFQp6KJ0/UjVPTDBh4ADRz0Ht5pl1Z7xM0AEAQiss0TXdFPEAwUq7wCIRmKbJ9EbhmYvi0HkP3df+3PAWN5Myj6eJbZwbdcQi842Da1DwU73CLoHwsMG+RfOqlL26mtmaZy/ZmP/DbYjlqRUXNSIEzL0FNZghCpazIPcYBDsj5czw73T/uQW1+Ok3eBtCGS15j/rqu6ApSRLX/I8DnocqZfjA2ABR/pep14L61rwdLjenuktjruaLbini2lOTIL/YYsM8nklXmTwfCfT7sg88P9U+Qt5Xi/Xj/y0W5+GUh7XAMeeVWP+Jfx5/vQQ4Mu/WldzRiNP30jK/L83cmsxaf1bJW92q3P6xk4Iq94td0OBwhjXlztSIovzLKTn0Aq7M9Fmf0mU/mw5FP0n/UuPp7+ZNzwbJmkduUXOuSsRQ/OQ84ToLG2vnjx4nB/93gSLE/pdLSqze/pgemBZx6YANkzh8zq9MD0wPTA9MD0wPTA9MD0wA/iAXZ3JTysyI1btgGZOfYTAtwbNTAoJGhc00ZsSQCYgLvIExyPCNIMmQogK9gNODECSoPODvGl8aPYfBLwVjC/7GvrHVvtrUsFqs3Dq8WYU37WHdOlA/ju82rpcX21LX0L/RzbRTq3z3Umj7T5QGCf5xJZBG7UxcBYPaQpGWVz84ysMdZxnbGziNXPgEfTFq/hKweNIv+W4xWpq4eHp4AYggDKVKf4ogdRV5YAgaVl0EAFewA10gZdFa64o0bREpslRR5g1/r6KvTZbjv8ZJ/gReZDcMyiT2XJeDCE3Hu7BxzTd3YfzLbh/pqMo59+9SaZZAEwwdhiy5jfs85hd1lX5W8aRyn/1DqyKf3az6fXV9N2f2c0dV1gtd/K2LSdXWddXj0P6Uf/rtvHP01Cnr2CON5f1mnG8NV8KhOPMbrrE941RgDK8b3Omldsg0/b1Vf91rRZB/D06scx2R4IP1WKPEEn9aaBVzKWrjz/rg/BpWzPpP/p6Snj9+PtCfJTptsLm7caK1vw1rPNlGfd4jV65Awv+LrM4IEgblg7AKKuZ33WZ5ipl0UwU/q2ce3bVMf4OtgfOThQaMwXCxx56YO8sZxx8C4ufI+14XZifcFHnrEfWS5TmtIn4Jc+dZPWDDLyXZq380UlwJq+8a2dTyBuL168XF3fvoxEbfE/NcwyPTA98HkPTIDs836ZrdMD0wPTA9MD0wPTA9MD0wM/gAcICokFRUY2W85Cf3v34eFLxO72+8cEk3tjf9MlCBUNaI2TDSpz5pbRIyVb0AwYyagQjDGAPgfIBIwGpB3YSi+MYzBage8AbxgnTYLYAdwIsITMQZQaswANoot85GdsOgJ45ZmxEb1rnLz77KcB14SnX/bJu3X02vchcrtXdKuMpNg2aGxHy9INHmpDE2W0pX7h33wzbmGc8js41x6ZyE26C62M+fAvwIBkjsNPAgqYncwgg3NBgjhFVfQLaIJ/z0vrY/tp+OtMY2YM8xddBC70q9li3ppG47JxHOCDGWKHp0e6AGN4m6G+Dm8dIpIRe/AfmUusJNoECYY+9CVbycwyfYLMV69erN5+8YYkOXgGeaizogRaljornwHnb8U5PiAM7GvNpDXjHDtMSV/zKjoBI8YCEOpf6fZuO3T4UFXw6rg4B0vgrGZdPxTglIyngDOCKBaAmWQQlR7JaNQmqpEzmLeIolLmAETxX1SQJ/b7aZCp9I4QuBTwon/bLnu8l851a+mthSqQNvSuNVT9zqd6cZjWasu9411bzrdjQczTL1BnnyBaClfHHR5PA1BkHP2WzjYNKCZgxidnmfmbMuxpm3xDrRyd69iHj6MDvKQJT32ScdiAX06AYGpvHxqkryQzn9itnZ7t53OQN2/yvAi++XGMvJL1N+YiIJvrPfoDkLLufUuodP7GWRi5eqJd8Fw6Zid+AjBfPz7UGzivbq6Px8369Ge//MUYkwtfajv81k3zOj0wPTC3WM41MD0wPTA9MD0wPTA9MD0wPfCjeCBxOIHdiPbW13/n13/xE04c+wkZIddrwS4CwOPTE8kyO+JCA8gRgBskEgjb1kU2feC1wXazlSZvJqQ/94oz8OQvUT8MOmMnXXwlWKd9yV851hO4M/bcF/ClAuMzTcsadPJv2T2u645ped6rd+vuNWAYikrf26Sah/QJ2P8/xLntr+bdsrzqxmovwML7JZ3y/JTtjihf1DiFV7+6ngjWHzh/7OHhAcwKMCfATPPX5wjzc+Zx4dt2Kdv785ZHaKNPrZSMPX+5DpxS5QAumenjWyeBMuABZKBO0ESm4912akaPDFSDcZGLPGlZb7Q9rb784uvVi9ub1WZ/j91kqaETjMMrug0dZdP6ev+8xO+F+6TLsZpvO5Jrfm1YlNAAFh49o4u+Xp/uI17Oy9gJm5G2m5HnHGT9w1KuNPlNZYBP2mB9UZRhWfJ+XrfPUV4bSGr6rNHoWXyVaV/zlVcX7c46oV+QpmjazrLPZ9/xTulmc82acl7hB2C3251WV1c1z0+cTeZvxAY/ZatnwFPAJAba7roo0FpgTaBNYI+eTWVzmSWo/H5jZtuxuSr5AmjKtd0irb9BrKyq0wz6RH/ZLVnbrUsPK7Y5DvCqX5RxCjCr5QVqNV+v8SvO0xbHNRAWG2F+ACyVJtuGs37QjXHlTwAx7N6wxdIpFzzcHx/oXK++effd6eMd966BUlVxs0wPTA98xgMzg+wzTplN0wPTA9MD0wPTA9MD0wPTAz+IBxLDD0lXr16/fctGyrfbze7qidSxAF6k0whwGZx2cC2924cugX4BNAIiBqhdOlg1UoYiPGwrYIG6QbeRbAe83Nrf4/oqP+8NLhMsiwCYvWR0OkoyXMa9Aa31jKHNgNo/MjkS/BrgJtg24ObTAIiae44Qjef+klt6lq7Fd3k/1IePQ4df1K0zrM52Vv8GoKEKmtLXQIv3NV4d+Bej9HKdhdUyHet9IB4Ge191/M/AR8CIR7e9CUZBe+Fb47RTX9ZZTA2OKHvQCh6IjpRBtDsn7auMllH1QxParQyFBtSbW7sBGsy6OWlv5FW/9sg74JkaMyDnmHUbtF9++YZMAtoBJeQX27VZW5XhPSBF2mVOqS119DKHsTmtgigFChXtpT66AyRK3+XMl/Wiqhb7/Zjl5zlV3u9Nr8TH5DRlXVamG8TOe6mRK6SfFGfpLE9eEKtbf87EAFO2xX/hV+NavzMPBizvHV+gTenVfV4FeBxvQfVkyNkWGuYPcfVoCQSR6Gf7aZzJJ6hU5/xV+xawrLZZstUSYOi0r2wwIaIAZqwht196L+jl1Yy7o1tqmSP1aJ3UxzY/6wfPMkMRSgCp0W79ijl5iC/svwCc0jtWeovDfZaTMUbFZyn+Hbz2gHtZWOO3TT3Sz1wVxIUf4BO/wMtr/MGC8PfEpSH4J4hmFpkgn5l0eU4gv7q6Wj1+s1/dfXzYmMF2f092pM+VQvL81xyo6yzTA9MDFw9MgOzii3k3PTA9MD0wPTA9MD0wPTA98MN5wAhzWXYEdW8IWt8QyO0Oh8cEm8mmIPpLoAh1B4wONCCt9go+bRP0MLS0PbEgVwEFg8oOzENnBLsoTV9jChho/s1HGnlsjU4p3e69fQnKF0CO45el5TuuxzquM8jkantnjix1qjElx/vnpfg9b6169RVKIs8lXylkV7YadGM7f5aMACSpmzTlq/1ipfQiC4cDzU9E8Ibh33zzDmDCuxp69oMZLKNEJ+6F0JIYiEj1suQaH9X8VrtAjmX4Lvd8oe+KN1mCjlBBB0ECgBAghOAAsdXD6+FtBtKJ7LCyq4DErBeyziAIx2zXRKG3X7zmHDK2xY3tjPa7DbN189p+SBujW8Mzr9b4j6yXpo/PY2/Z1j6Vv+a5jHbKH5lUKhoar6gtH7fn2Z925KkT/1K00XZLtdez0esxHePL/qa1SZoGdM9AbjOmv+n76pge77Xb28aAVehju+u8nldHMU5DLQv+8tgMUE2ArHhrG8ZpPEXwS/4n1oHbR53ZyGO+j0/7AEiCRw3OHQAWHd+fJ8+xQ86WNtdtz6tX6+olMGn9EXmCUQ3q2bZjK6jAne2hF7RkrR/JLPN3JzpCpwwzyYIM0mgmozb4iDU/aTwrzS2VbvHEqoy3PTYFDh12wzN+CIX+q+f4Ab6PZHF+89371bsPH9dvX32Bsepxfv5KqTFuXqYHpgcuHpgA2cUX8256YHpgemB6YHpgemB6YHrgh/XAMlDbvnv3zcvXO0+TPm53BJtPbikiMjTINCQ0UK6AcASNBJaCOQke6TcTSLjAfwa1HQAb4Pc2y5i3lJoGQQGDywpCDXrlWUHlkGUgS+BrXG6L/R2cVuCqjgSg8k4mTI2TvUG7JTzHtcfa7n31mR1Uetje5UJbil/oayzaRixMSid1BzDxnDaLGWLyV88E9GTkROfqZkwDihcAIoALuoQFEbxvqzRgt5ySWwVf05to2mxvw9/5OUDz23/516uHuztif7NpDPIvwId6+CeQ5RypRwEG1BtcpE0bzb7hRhFl15kN7TY6ltWhRmkw64ztc6bXbLZX8WV8Z7c0ABZAG/FNtl3KBBnHg/PG2jpW5pAJNj99+xYX7ld7Du3vbXK1XW+AUI4b2XNyt5SvEMN95lP9Ryk9lIMOqoIfYqP2mUUkqDXGOUcFttZ4rMLTylXmaNNtAn4AeDmjj+dFmdp1gFfuqes/S+QLoiFFfrpvDRDjeHURpdE3rZNj2iC3BZqdGQXTgT5mZY3nJLxDX+vHrZ6xXxbaB/+uS3Y41lsoXXfqc84OPGcj9nrkyY8N2Ip85bV+kcl8RgdALDNKj5zddgV9QDKu7nw8CJ4xVn0tAli8DCRXPRPd0uNyGnrLY9BHpsCoelBK/obfpqL1zLhHssEEuMDiWHd8nspe2zwX0asocOu/5Y2rfU8HtsHXSXEBuTj0tc72Vrn2O4/Ot42sMOv6RN5u+wx4eZX5k+D07YePq79992717uPH9e3NqxzZl0lnOuifZXpgeuCPeGACZH/EMbN5emB6YHpgemB6YHpgemB64Hv1wPNAzf9f+ppzf14T93noGEGkAWIFdN4btHbA6LW3XqqlwXDiS9sNyq3T7r2ZKoJsxp0JNBcxovWc2STdAGbkl2JsqgIwozvyDUgd4ye6QGif0qwH8KFW44YuoQmRhCnL8d3mWANnI+Jl/4VXU7Ydz+rI7yIfgRdLZ/50n1f7PVtrKcf79HFJdk8CdYNvGnTo0Msg3TZBA3X2s+ZNgKCaHJB+WL0jMD+6hSxAjQAWJTxKv8hEfviKRmWy5Fl2BbBxiDOIjIBp2ua9avDl9tgAUgAMGc62ztX2eszsADiiv7AlY4e88JQvJRlL6i5v/cXcHp84Ow2GV4AN8t2ydU8cUF0L1Cj5jo8djL3Mz2VN2G/JnA6aotcMfdL8SpcQjy/lZP5QQNUs8RVXZUUXQRJtD0GtcYSd+3udBijWdYphPgROLQF89KPAoOgMzoy70nv5Knk1x2W/81S6S5W5byWpt572ee94aT4pqBEA6tm4gHBnmy685FF2fsIl82qWlnpZztcht3XR21vWRuvx8uXL3Js5ZjEz0L72meOu2aLYuvfVdmW49bvvW6+WtT4AM6KO9S0g7Zatv9Jb5G8xm81xnZUmEMzTKEZZNNaRI12ujh/rwHqBpGWzersSGtxXri2PoHUCdwDF67sHz9FDsP7+w+UWnebX9MD0QHlgAmRzJUwPTA9MD0wPTA9MD0wPTA/8oB4wOBwB5Qj7In63u7l+Q9T4huB9dyB7x3je2Njw329CbT6OFTwze6IykAhXE3DKTL6Dt5UE0YIi0mwSp8u06Dq47eizxhHgKtRgEpmW5pcAGh7yiw3QdNAtHS+Lo8ecmLN9Nqe0zV7VRR0Ml607wnttWhZBoDNYFLuq14PwLb69M3y5T+Bs+pn3gk4Rgd1Exq1vOvkSGLO0XanwZYZcABTlootnGzUNOS8MCNSUPttPe4wwPHeiRtld365+/+27tBfooqGl74mMwNKwiG0VqKlsLmuZIPhBJZAjcQM6yKsoHx3ip6JVhtsmUYp++JOdc9YG3mZmddYVzorfizG86TPD58TB/AKCAkUbQL4ddr56cZPzxw6epZblpz7MboMWZF5tAZesC6g5D/rMq2Is+sh6GtKuDHjYr218Fb0gFTUQErOvely26dEm38xvfOHqcqSZYwUEnuxXDO1+1Nez0xxjS+bKZteCgiwBXapPOfSe5Z5pQshXmDq+tiLaHLtGv/c9prLB0G/IWT4fg5y+skmajB383LpsVp7FrDjfDNlgUPlpPJeDPnTYmrdOhnasicwHvw+kc7WeG2S5+gRxPVNNva6vOZcMXfQVD8pZZ/mqRvkLoAoat+f6sai3H0ElxMlOAAAgAElEQVQ+z/dSxsEsNp8RytGUMApUgGMc1G+WlzTqSFfPp8uc0egEIMcLA0Ln+JhRtjKs5MkP+mzhZN35YgAP5Y9fEKtNAd44X80z0j7c362ekG2m25GXGtgX4bFh+EklZ5kemB74xAMTIPvEHbMyPTA9MD0wPTA9MD0wPTA98H17oINn5FQkWQJJHrt+zV6g1wSmnG99CUaNQQ2UO9iV3OCVEDLgzJJJsaqgcnnv2BF7J+Bs/ra3PrZVUHyRVX3WK3OsXgQwOFckG6DOYDVjVYZANoGr0S0lTUS3rf85s6sV76u0PUa9+MhTV6jHxv1blHNgPGil8dPulLbtik0E+JZuk674ja1nQ35k6VVlG42PMYJ01p2DbrdP3ue6CA1FEOC77z6oMDXHIFskwCKNYMPQuxovNjukZDu33FMfI6udcZnz1s1sPpkIknAjyKXcZJxxK4BYgA0O1AYBjPhJ5sOmMUY22fIpIAYo9QKALCk98HZM+sKPurSOP6/JatMXtj+3T/ru896ypGkfCnjZXnM56GDtk1D0xV8gRaAk46D/tOhfR1RpmqX8lieFfKsej1Nftg0mXJY0zoo6tg25B+IV3FPbz2Usyql1uMi88LXvAMBpCTjmPGK7tL3uvF8+t867bUKia0AmeUQGfmx+XncC6Vwd60dLnTHPl9tix5YzxJKditukP7KGvfrJof7DVte2dIJTriuGD/0GuKbzKGKPdX2MPPnE5jG/kQHPnS8fYK3x5l5+m46rJ+h2zG1vJVfXfjMpEhQWPtxEt5JSWWfhz3ifsUe2Bd/x+cCbK10nr1+8XJ8z9lC9x83r9MD0wB96YAJkf+iT2TI9MD0wPTA9MD0wPTA9MD3w/XugosmWw4FI+8Pxlo1NtwBBmxOBnaGvkSiFJBnBqwo0uU0RQDIwNC4NBJTQz84RoRILGowaNNaWQWip2nYOWrmXh0F+gmfu3a5km6F0MosAHHoMIXL1oUSyi5CsbEEBYmZuolp9wTvnco3A30aDecwLPxWX7wXOKN0a4Ihe6hfGpWP0to0/RWV8GFCDn8VgOudAhS5N+SqcCq8ShGsvVMm+yVsRGSpwlz+Df/WCZYOKMhC4UIL2JuDmqs+cD3n6xsjv3n1YffN7MsiClZRvlaMt8o6OXPSjlhf4JlOAB/UPiX5nDM0owhhvqqhXgCuquWWukoVmpeXkLDLnA4mso9XuKnzDHz31Xd6GiI5m6VWmlmAhMiMf0AS+Uu6xzZWg3AZ+HJPVAY1lzfY9+0eiXNr0S7L3aA/NmBvbS09lu76pbSrby3l2zZ3MavNssPhWndCF8XmDJkCKssqfsFIuY1rvIS5ulqaLvJIpBUH+uJYuUAw6s6FcF+3HrD/qSz5a43xaut0DrjyLq6Qxr8rgk+2dXuFvPTq47qDNeLOy0lcyylNIPx+iL1+1qbHOm3wsAeXozPmCtrF2XYOuyz3bC0tWnQ2WDDDmaqefGNN6V+ackF7xbT29ykdZHpbvc+5qVeaRDMV+k+aRZSXd5sRNdKo6T1Xq5zbWcp4P5OT3xOcIu/jFiy7mcyrLl0IcXR/D5+rRbyY9kg12BqqhlV792xa95JbOAw8DANn6/cf71T0gGTpvsOEaFLB1qins2rxOD0wPfOKB85PySeusTA9MD0wPTA9MD0wPTA9MD0wPfP8euETwQGBsz7tl++ALtvoRq2/cYWWQTfRqAFtBrwGhW9q6GCjSTRuBJfcGitIEsBqBZFMb4Bo4G6xaOshOZdS7zzb5EpUOvhXEdkCqXAPWI0G+YEYX29EmVWkDJFU1bQULXfqLvkcX6KBelgYGagti0Szle++ngRs0rHHoYLu2pox6+afstr3G1pi4NLwKCGje8mwd+ypXt/VZl06IwY9af8eb8+7IXEF4PqEZLilaiAQwSyw8CoiQS9vtlrkugix6Ylmi9/BRt+fNlQJ8ABYBZugXVPKlAdpt9t1R4IwikBVb0KHPN3Ou9dcJcGbNuVEvb66hLNClAZEMXny1/eEV4Kr1dk7Kb+ljTM9F1atP1WJL1hDKxJflh/JVOcmx7Rszl6In/C3hO+4xHBY9J+kO/5JRIFMDP/aqS/dZFyDUZhQZ19KPyig1F8txpWf3X67Nt+235zxuASB1f/e1ndI/522fbdr8vO/sE59t7BKcrOez1hrpqVglOOzcaF9lcFV2Y/FrXVqGOuzgc9y5RbGyx3xZgnpIK2B/hC8PwwDUCnw2CdH+/sjHkt8Crm0H3g+4qW4+B8ol1Su019eV1eZUyCf2aUr41tU+weJaEwW+HZn/+/1p/fGeZ1BgeH/YHU/rN4CEGOmDlDS/WjyRNL+mB6YHlh6YANnSG/N+emB6YHpgemB6YHpgemB64AfwwHPQg/9LCib2uD9w8NOB87F366enp+MTh0wTEK53V9eE1AS4CQYNCAsYMNBM4EigagqNwaMlZ3NxTbaGTbQnoPbeoLbRGWkJSpuP9wlAabd4320ZL4BihziCwekote2S4F16Ql40SU99l4zIcZDyB1/lWsLbUQzw/gwAQBvgJraVQMPb3nYlrVuoBPVK17Bb7cQUYdZ6ROswr36zwkIP/8ir5oTOggjKLJ3oYJwYpeeRJQNLWvQ0a+mUrJQCCwz+1+vr1UfAsY8fP8oARYnoQaM4Ui4eyVllC5udCTuUhRRuyh9ucaOCHl6546K+oFfwq/ClspOgkZ/jOFsqtPIKLeLtAxjbAkAUODaAkPDVCfbrnfIzLZLnHZ03nk+FTcvtduoUvzhGv0QiX5zNlTkTTF2U+GvoU3rW+NirjqOojh/BDf/kpe7SRd6C1lFKdg1Y7Mr6c1VTYcgoY2xXuWbdo6Nb+rrEV6OSs9+8d93B162EFnXoZ6RkOL70a5/YLnWeR+9lgJ71bAwQlG3KsWn40RHWzfCyuGW1znWrbCmfE4tbT3NdpujZ3v7hvvVyNs3adM0WIlT+DHAInecE2u9Y3/Kqz7239BZmpQZEQz7gErZLu1pdsTL6mfWtrgKKsVs68KfMC+0uO9eOYHiDYr0dV5MOgsLYCoSLfOd6n5dCSPukXujuds5+gUL0c6D2sjbWgLhmlq3hw+rO2tHXjkPf9SNfT+gckHC7ueL2JzwDX6Hs72BSCFwsZiIwtW7n9/TA9IAemADZXAfTA9MD0wPTA9MD0wPTA9MDP4IHApIRoHk1Ttusv3j9Znu3P2wFfQj2CPUC1SSANUjcc5h6g0cGph2Mq7z9th3YisQBZgShFeTb3kFt03jt0kCE12X2WMbAB6ZnYKhldkxp3eK1PgS38FZ2F3l6jpG6Zgtfglh4DprSSbChbHCcgfIVb9Gz2O+fMo+8IW9Z1HHpA3VY2iat9bYtNtHWdOrqvaXaCvjp+qd9rYe0Rd/yncM9Af2ONz5+8+7bwVNdC0LyLYG+5ZKIvQYPW+XfMsoPUWRhA/oBI1jSX046jym34EtYFxXskcFuXcA1rgB0AgqH/VPa9JU6F1gFUwGXgEG1lgTSDo9sewMN2ZFplLls2eh6Ht96q8+5FDDSdtT1sg4ka3tdVl3afvVKFmR3jKt8GLnwSfERPFm+bMGxvrTiImMhBA7yie1Onhy5Fu9Uc9+6KLHoC9hyDVvvMXLoM/nUjY5BL2hU+EuNr/Yep6Tl/bLe7T7xaeer21Ifeqdz+N1+S9uBhcydzx9gVrapArgxl85b0ehjtlry0V/eBwg7A2/ls2ov3voMx2olYDTjeS61cavsHb9JPNvtV6+HbMGs3xL79J30/gm25jw1gVDG2+7ZYydBXMb5eG/g8chvmGAyXvdnMZ+AmsNuL453q3aKNJTy13b1/sPd6iPbK5/gxe/MFY/Ea+x8A8k3fJygGsDNLNMD0wOfemACZJ/6Y9amB6YHpgemB6YHpgemB6YHvncPNJxhgFef1z/5KWAFqRGkO3hWEhlkq+tsPbKJwNSAkEDXj6WD2FwJ98yOIVTNmxjBPKTgQ1swtgpwE+XSHjqD5LG1jTCeOLT4miliBNnZJHKSjyUUBJ2VFVNtBqX9idxRzwBGQM7ozgi5xKUGwI6zV8AmQTwCqAXgS19kCRKVjALKyvYE7ozW/i7tk+LbrXUN/UAfmh9sU3B5gKQzcERHeOGIAHzj7YXaF1sdxZieDzOAtusCDr799ruAAPnv8M6bfmXOopP2ygQnJzsI/yc1J46Tx8iMAkBIGlvENJCRWanxzh2fZJgBFHU5qacZZgJxvLLUFeF2yXjVeQGQSAbO0Cdi0F0/yE87Nlc7cI+n1S1Ziw32xGac1NsXXYsYFPfpA88G8+PayfrknvP0gm2om2tQ/lgS8E0+8ow8dekppC12yf8zxT5Xg1dXaV0vhPK0rdZuMbXe7VIGzBmPnwCLmXWhka/rb/DQPidZfzmmZKm3XNQiLki76tR6bIAV30Mo+FQ+1P7qk492a4n+tzzPqIzchWzUKvmsk+g69HQnrrJ7i7F9fq7GklBX+9VWsFNQzyIAarYVI9Pu1SJN5o97s7/kZfZY2SIt42m7Buxte7XFezPKvCrT+TR50nJ/f796FKjF/kfWo7JqKyt3jA2AhiMe+L27ARKz6PMn/iPBSWDS36jMl14oPWMGt+qozlvBQK6Cg667x8Nh/cA5bPTCnw4fRol0Bc8kHcWIhlmmB6YHPvXABMg+9cesTQ9MD0wPTA9MD0wPTA9MD/xwHiBQM4Ldrf7Nf/CXCRZPD4/gNAkcDezS9mhGGfcGgwarFgNZ74VBluFegtkBAKyNCaHpMXWlMzFj2CQI7mhRuUSQCVClNUC29L1176XrYpBafEun7iv9iqr59La4pR1S2N+8O0C33jaWgQJFAhFGt61x6XahK16tT19bfl8FwlpeoRQCAQJUZd+5D93kUePKbu+7v3VlF1eAEPGub969QztuQmeoUWCJdkZtjWj9K1iHtOxRh9LZOp+BHG3ITAt4J5Bm1oxX+aCbdBnDdjMQhdAJ9ISGs6PMstpweLmkslPnI1s1a0xGrzYAHge28+4Ax05P2AvQcANA1udC1Va/8lH5Av6jxD/Qx39kAnltv0gSf7mm0NdtdVEkdW8dJ80ASOObGhO+1DN+XOW7ZoecHgw/jFrSeS9Ntynfewd4VbeMi/8L+JLGUvwu67rb0slXjy260guujoT3ct5qRNHVfcuuWoZEn952qL+j5yBwbJdqr36fG4tt+Yz79rfj/BT4pU7+fni+V/klg/G1oFSX5ViBqKYVVw3oBL/dAPcOQ0+tloe0nKrPvZ/KCKvsUeaVuiCZZ4lZBPylf8h813rRp5bwYQ0+7ll3yHNr+XY71sRiPYUuI+qr/SQIWeeY+VKB0+qbb7873ZMJqW1P7LMEvCWZ7EgaJcxUPiti3BWr+T09MD0wPDABsrkUpgemB6YHpgemB6YHpgemB34UDxjungAv/uE/+ser//q/+W+zI87teAaCxnHEigFekrFDpQNCgQ4zN6QyCNyzhS5ZUCP4dFx4nONBQIOkhsGVvgKoEg3H7uJb/A1ZxVe6GMSaMSK/Oo+KmBgejukAV1p1qsP64WODGUdeR7vjk4FCE7fp6EyiDciSW6gwJVsE+zwtdVGOWSSWRLcBf6rdttjpmUYwzVlfypFP6jXuQldgVwEI8Eg3dpRC+BTbMcSxTkBs5D5+homZLWd5ZsiMSMI2A/R75u79+4+R7xlKMIAhRIBUVFSqeNQEhX8f0q+OAy1ygtIXkIvmyERZXt6Q+wAq0uAzQaY+q6wyxwTKBDrxHgiF66PtcJxzlvHy1UiK/dleeXeXM7CuSUG6veZ9qvDfY1PPc96sCVvHO6aLb/8URLFUu0BUKvEtGgYcq77SoYCZT8EaV540/VIA72tMWJ/10B/JZsNG5VArAlKLzFbrdxycx2OmNtTcCZTVGvEaGkaXX8q/SYUrjvlmZXItX9mQt1CqW3ovPmx+yrG4zsJ3AEzOn+diOT/aLwB1MLsKnaPHENHzAuQEuFnrMfqPuVyztjLeeY4Dyo7yi1pVuzS1/RY9oBUATkbjsNt15hhBrfaVV+VLf0VGFyzyXFSWm/Mr9yEvD4w2xtycI7YLL7ZV629wOM88M7PxdPJMO9bJFfICXtW4yHdLpbbwqHC0PnIrUzb02jx8UBlwOmn8RrI+d2aZlXj8ueXNlY+cA8j2SrJwBb/fvLjmPRXrO57PO34E1bQW6nJCx/h5mR6YHrg8INMX0wPTA9MD0wPTA9MD0wPTA9MDP7wHACD+w//4r1Zf/vTr3cP+cE3oS8pFAlcjQeLHBKNgZBU9dyDbitY5PlWTxkA6wXTTF5MEwvYXnwpwm4f0f6yYKfKEjga8CZ4JqpclMg2ph7xlX+gBr57rvKRZ3qtHjSl+3nf5HP/u87qk1SdN79VP9+OhDEs/Afz5YPbBjJg7RXo/4oomeDW/M58BLli3Lz5n8Pv371Pvg9AH2/NF0CM8zB4bujTC4JguyRgbFfCTs/42WUdI6dQ+UsnQ2a79+BIa6eJXYIElT/kEpBqgDevOJkCxw+qarKOyqwC2dNjXPhE1GfX2S9djW3oVffH7sr3v22+Se98f69GNa8v0aluPlabv+9rjsTql61akaTrryzUvnX1euzTt82vT9FX6vm/a1t0+2/ojXdYJV88Z9L7r6ROYGs9S8+yrPJbj89w/H089NGO9uJVyCX6V/wpci07DXO+7ON6Pba2bfW1Txg368KPPN2MKooOqcS+otmGb5zZtvHAkWWS3N1crX/xww5slBWBLl5IhT2XqE+3y+sh5ZwJk/ocA65bWzXvHLHWqto0vyTh99+Hjicyx+JJsNMw4PvC5l4aisW3wZcLTNb+mB6YHZgbZXAPTA9MD0wPTA9MD0wPTA9MDP4oHiM6I8tar+6d7Mh8eAMieXhDQ3iYIBarYP/JONwJBs5MqpHNbmEEjB/GP88lU3AweS59lZODYwa3jBWKCx3BvlpUZOjY7Kv1UDMwDBnFvRpLjk9mVMR76L6AzQBnvRiDN7TmgNmtMYCbM4eFfAnQFJZWl9HSMckuPC3Ah8BPwRwILOkhnpk10Xcis7gK7PHNKfbpss6Ww6mV/9ZjkJFloccjxINCjfL7lrRwJojtd3tqpUvo446Xbkrkysp0gEjMU3Prw3YfV73//DWPQh+H6MO9ZkAC+aw41l32+vNJcn+LvGwXDLDSQIW+pP9SjQKAx8nViQ68+zCLZOB6kLmvPsovSnCkWoq3bJsnWEQU0zQoeemDjWnrghCjACQGKHSBGvwk0vtA3Ko4PFOU2z6IrIK3ehEg78l1Dli1rEIwCH1SDazLZRPph+JmNeVCOtaefGVzbcAdwov1I7C2oyjRjrgy2z3l3vekrHiVuCnghOyvjam0d4gdodJU6dUZXBqIrtL19Ud0v+skY/dVtUc4ZjfSVPMnKrvNY9InP4O08ZXspvlBHXSLbgJjwrszMWuu+zCHrRpkSUXyhRfj6lHJPTl+AKB6uM0gknT4vPThQH0P7+YUD44t/WYtJxTpXfZy1j39jD7yU1584TQHSqffws750e6X6WjKWftTIfNjm+3dXR7d5kpEGMOZv1M3JF3C45RLw/QkgTKYUM+7q9wK7PEvMF07C7AqfaE+epVAO/fQldYFAsxqfWPvvP95xntkjgD4dfJ2u/G8Lp0c+brHMv5gw+MzL9MD0wKce8H8TZpkemB6YHpgemB6YHpgemB6YHvihPVBRN9k+Zl1wSPUVgeYrAlVOjkrgy20F2Qa9lr4aiBZYYMBqX7GS3mLA2rRez4Euwarjqgzxo982af00qNHj9gBqaUcvdXteWm5kGR1TwovAVV03AC5dpE3fM7m2S2tZ3j+ntc/P5+i6PZ3jy/GWvkojxJA22Ii3JNMqLZ/ShSb+KABAHs6VRT/ql9ZH0Onu7n714eN9eOassCE7Vg29Iz9bLpHF+O4L0+XXoDfrq32w7Kbxk6p1aXsbqGePtW4iMnhNgXwcVmtCQMy14ttRYxtA2eHAYelk+lxdl522L+dFno6xbdmHsOhjW9lY9bMO9DpuWXotNa9et45ZlubReijDTwrAyLLYvpRjvbOamo/9LaOv8miefW365v+5+nLcks77pm9+tim79bPdT9fFLfu5brq+dsZZjenD/4tfj/EqvcBkH55/4c98BcCu+Qm4utBR3fSvOjumi/e2WbrfunK6XQBT8LPnJ7SuuDFOYOyWNeW2XdeW9G7J9aUUjml5nUEmb8Eu7fHjvW0lv3zWvKMYX/SyzNer7969X30LUO0YNPY8swNnMYK78UObom2frsNqn9/TA9MDemBmkM11MD0wPTA9MD0wPTA9MD0wPfBjeIBwTvBju7rZvuBcntMNSNILssY6aOZ4sl0i1QSjathB6FHwgi4DWeO+cTtwstiSTB7AA8daDL6P0Ob8KZo62yzBLiwEEQg9SwYXbqruXeqIGUGxdI7rM7EG3uTo0omL8ioOpZWIPSH2CJg7uO236mlDtv9B1H0GzacBmG1RwGyzAx5L/yKAV2QAIMScyKgJEJTGCy+r0VcaZFQgr+/LN/2GQXqhgxi62Ax65VsO+8wys1sM2OWlCnVVN7aY3V6tviU4//DhjvbkJJWwoYsDkkWkLg0uhY9KyQxhAbC8j8KpGuRrU/xhBgxzegotumYoNgw/KepktpRHLY1z48LbDotynBSBEujytkd0OLKFTfxAwEzfvHz5ki1yhElHToTSYZT4L3elpvV+2ULOJKPPjCV1jxiuqDu+uCraS2wdPKkH+OCgd1t6nXkuVwMnobcPefURjEF/x9qekTX2AIMrfFPnkxU9JJEd/yHbq3y8bsimbNyk5eSKf0KjOQjqc7vKNiWX/r1+IsPWwbev8vIjENj3CF1t8anraLi2nhVo2n75ycO5r2e/nOf6duNgimuIAemHVtxWL/oChgKSGJ+XNAAQ8hIJnx+fQvnCNVe96HMnPaamyC+/BeoObdHTNe7VRP/7JkqXXfwV++Qu4IXc/PhgD7Q7MhX3rjVqrimOIlsdb3i7JRlke0BcZflclX9gqHmP/kcDfpPIINtzcP+aDNGcQ0ZdurN/h650pv3+8bj67uPd2kP+j6z/x4f96uXNCzme2GjppHM7y/TA9MC/ygMTIPtXeWf2TQ9MD0wPTA9MD0wPTA9MD3yfHiBi26x+9rOfEwgeb8ncqu2VFYyaQZaIzqAwQAIRKXEucV4FyRVUEkASoC6L8alvsMx2JXgJhklhYGl5frWtA22zTAxGz/VFUOm4HttjSoeWX/zNnsqWRcZKL41BePN0rKXrBtw1svg0T68tL7IHlWO7PXywTh5dHGfp67l9kKiL5cAWrAT70HuAuX5KT5xV40uOAF7Z3roprvl4NdB/eOBwcIAPt78+sHUsCAK6yddy0edSF/TAGHr1QSnYwIljlN/jLveMgWfqGRvmfjlk9AnSVQmd4OaV2TqjHyFti/qLs16xNZPX/a1e3r4A3IK/w4d850qQo0rr1NfRzEWe4ad+o658i30XG8q2scTT71fksHaXNtdwFBwWtd6xZYyUr8e1l4xq9F5dlO7VEmAKH7QeDRjLu/WUrmSUxMDRsaeyHM2wlPYCrDqida+MqIuOPns9E0Xnt+ulMxARlg7HWFo3pZsJuB1biKsfcEqAi/lYFv3m8BMgpfc73ny6542kmYtNZROyhPldAACDZhMQaymruLWfmndkxlYGuzdUHghSf/WrufG+7Nc3nDAW28rl5attthcDkvFs3D/VFnHerQoYps5suCTjq/QvfzlP4+gxXiBRzx4QedkDYeZ1zKmy3Sb8uL9bvQegxhO4h/VKG/qDV2+2XEtJiWeZHpge+KMemADZH3XN7JgemB6YHpgemB6YHpgemB74Hj2QeFD+BqEEfK+4vUlAOtrsM9CrYJzgX3DMdC2iUoPFPuvK0H9AYA6Bn5AALQNpMWOpgnxBhqb1pupmtSTSrWiXcbX1qQP1vgZ4Y5iBdkqDKFRK7+pAZdgBTJBCZLuZKDnDjG71FJSyXb6W0HBl8xVAFNEyQE7bLHAlIGi9ARD5FSBQgXpAgPAbesDCIjRi9o5jhRMiRzraqh+vcGvWiy3lo+qTVjAgBX8ElIwu5Wnb5S+dL6r0+u23364efUPflhQZ5wmgMGlBysR5p4MOoH2AE2oSgEZZ0bD4oDB120qBShijjh6CaNovTSASJ0PFR1vGqK9Ze2xty4H9QUYY7lFkgpec0Wb2X/M3c0xJ+tTz27748k1ACVUQwDv7jXVUfmmfOpe0+YcN0Vg9mMPMcRiUnB6HGJjW+E/BMddKAVCSOGeOqXVQYJD3XdIXiRKzMkZf5GgN9W5zDtINmwBTvPVV29UXZ+ISdbSl5KTCV8vP3ENivfhf+pThGrMIZwvs5J52pKZHQEnf5jmj0yUun7zVtZTIGD1p8dt+z/fKm1mpZ71zjbw9Y1mze2is+/hm7liRB4AmbXSZCdQqVl7aX6AY3LHFhKoq8NJfFJ8jgHpoBwDGYPm3PiGiYr+2Rhdo+vnzWLtkkCG8z7BzvSoq9gL0+TtwzTZLIKtai2sQMp+/Bw7pR0/pWL4wBzRDFzZbrk73p9Xti2vkoQ/O83dAu5SRgoADPnn3/oMZZPLgEaEPenyx41m44k2a5q7ZVgu1Rs7v6YHpgWcemADZM4fM6vTA9MD0wPTA9MD0wPTA9MD37wECOOM4Ir4Epi8JrF8jlTdYXgpBbzIhDHQPZF1AmQBSigTfnUlGDV4JWC+j685A0vjf/i4G0x3UGkgmmKSzeSxpe4xX29NH4O5VHpWRU7zlW4Gp1AWOeffHSstZ8qrMlIu+9i31a16fa7PPdvWwqJUhtBFx7g32hx+ks816ywit8mh/Xoq+dOnD0NuP9l1d3ay++fY7/IHsoXNvGw2CIVgJcBA+3OaKnh4uT/oMGA+gxpiXHFQf1AMNn+us/n5oD6xi3bcAACAASURBVA/BNhEXwAcNck6SsQZNgB3RCbrWrBVfLuA4i6AY6FzuHRMUg35turm5CQAibbIPhz1tr3wd42fpP5mpUwGjzoEAT8nrvva1V31V813ztaRtvo7rMcW77O57+zXfImgTW5xvfcRMZmwDKaEqHb0t2uJvXVXlO9jZVPaNq/St41I/F0zkjJVTsh39qe0KkEdnjjVd+GIElvHU4BPojuqROXTNla6aZNtSb/W5gHKlv/N0GevWRnK1mDPBKbfBCpo6znUce+Hp1XFV6l450VEFKNJUKXrvW5dP+0RsnRfmQTlOjGAdSw7rVqTJsuQH+AaNeu0OrH+2UHp0WOuhR1y8DF09se1yc+0LS5z/wR99XT8t++P93WoP316n4wUCvOPgtKOtFns0O0+xApbTXb3ze3rgT9gDEyD7E578afr0wPTA9MD0wPTA9MD0wI/ggQRlBG0GZgnOCHBfEmi+SrYDzXcc9E5dBC3qeS5ZlQpM94Ab5zfxGXwadhIongPLGka7ogyWAU28tWZQSYAZkGMR8NpXWV8QnsfbWiVBqCkiFO8NjA3MvV+ze0ldk1kiT3Rq3aUTBUw/fL2asyJNZYSxfREAw3azjoqfPKrNa2QOnaTThtAN+hAsEkN665sBuvLPBsV2+Ao0BlUpf8pLnslg0jed+SZeoCpmf8GLrzTI0aw87bJ4lpXZLu/ek70C7xx6rxOhESDwrYf6pmwpmYJh8vB8tj5rjQHoIXM+iuKTTLBsTysd1FUPWtTTMSnqxrgAX2yv079mLoW3tg4y8bTYy1Uf1D3AifxiHxk+AKBRjawcd4Da7sdsMYtnoGVnqG0S4omohHzp4lqUcY3JP2Mg8KWEzo0gkO3Od89l+NRAdLVfWtcrVW5YJeFNJfwwDB1K/7MMu9KP0hR1sc+r5Q/ubUtPfXnIu38NIPnQhDdEZWfRLfnZIo+SUP2tD4zS57OXuYa/23qHG5PlFZ0EdaCt9c9aYTZiv1l+8Ql86JePWxjNnMp6hahkqUHZG5u5V1/v/ezXtcVyO3zXZ80dAMqk2+bNtoBUnsnGApFn5oixZmG1vWadlR/KWvWx+BxbssS994ayHVu1sz40mgXA0WDOPnzIIsvaqaw7XnTJFsneCgotPtFR2unh/fpDjCsfdOqxytnAlF+iPIOAjyxPbXdb9Bbg+trfxhMANkrBl3UDc4fNMj0wPfAZD0yA7DNOmU3TA9MD0wPTA9MD0wPTA9MD37sHjCL5HDdsi3rJ9SUHae8EnZIxxlXQy+BQKgNC49UGchIwJyw3oBdAICCEwNj0CMhjQJluguIE4YAVNiSwNPYMAUQBf6yXvfJoIKRaPv9deiAswbzX4un46AHDvq+AuQSULgSoDNGeBOPeEOCaZLUsytAHluJpcFtjis+QFV5lm2OWNKnw5UjtItzXiTKJbPnqY+X0IfpmcJV/kDsc03UBnpoLdaYE/Kqtab/79l2Ao7QLbIyzk4blNBeg2DhQQIAQP/saMpWTbDK6cz+2OwYE0meqIEg2gB1twiO02SEIICAw7MRmV4mZSSCbsZ+v+DX+gFZA40D/27dfwKWAEe3+xNfKQHb7w3u31en3pkNwStPYp/49vTWmQKCizOycx6i9peSoaunQ/Kq32i90Bd70GNt7XAN1raPtoStvSSn5J8V+S8kcfhoU9i3XwJnfwleDtHSAf+iZqlzxrQXys46RM/hWH51joezy7BdIVtsmy59b2AgcZk3KjzksG1vvupZPBJbLTg/OtxxYT8p1jalXeOUhdA0VwObcXnxRz1/XY0A41Vxlu+3w22gOf3n7eyVw5ZXTxrJs1wJbrMWbG95yO+Q8cnbfA4f6q8aRdDLBwD1ALRLyjK5FWflJuMZWafx47t8TdnzH+WPgj/UsIys27dkkfFpztF69Opbno4wvBXuptbrzOj3wJ++BCZD9yS+B6YDpgemB6YHpgemB6YHpgR/FAx2cbQkSbwnmPKB/Y4Br0EhZHwgWDXrdUWTWWDI97DIwNBDtK00eIk8smTa+CXorqPTebAr2GVUwbLZKCEfmx2gPO8aLrZC7FlpgCYdfSoAXeNOSgN4gleA6OhPACsjkzYhmb0R+6Vm6ZFDazZSR1lD1AAgQCEzZBusGwulHP67FJ53JptJIs7E8qFweFtUSJEAa8hkDuXrRmH5v5VPgkTyxYdiiTAEIKQXDQic4kLoDHTv0gM7+/QCDdtCteTPf7vpq9fHusPq//5+/wRfowRlXa/aFeX6U5cSbBX1rZFRMC19OKn76pIzsHTojJ2AeOsUvyLS9/I4lMaJsji9ZHxu30kkPpd15oyXZZDl2CVAkY5C55c9tbb7IIbyzrQ1dACTU8Rd/9jOyyHarO+bmVGux5MYXro3hWvyhIPlmzeg0inoLTuQevbcyPY91ncIgYzLzkKkbc592rNEAW6lHZ67yC0+3GtsOUOKYM00NSZ3e6JOxtNeW2PJ/Mux4BhQh2CJNZ/DJP2Ba8+Jqph8Wh2/uVJ2141sha9VoShme+ZJvQGdH6YN6lmQZu9D9ODIud+BCPjtmdHpFSOnPtYv2WY0Ps+b1L/Q6FPdd0RkbtElaU7QoeeYR2PNgXyngmq752PF2SwTze5ARjK/1jiIBsBgc0Li3ewIhF28NgR9mRmZwN/WwVzmfKTV/dCDCzLUGy17cmOFlFhtztvLsvsf4Ys/ceq7YI8/NFf7Z8ELfx0fOKwMa27J2tfnFNS/+VUfGP9w/ru4fH/LbKYh44mMfwDcSV0/bzY6FE8vQU4NtnmV6YHrguQcmQPbcI7M+PTA9MD0wPTA9MD0wPTA98H16oCPIijaDA609g+wlQR9YTYK6DphJuACQ8Y2IBK1+EzemSNeZTjnryj5DVINXLgatBrCWBN91m6ARWCCBbbbYESwaLyfDA/oE0tAm2EZmgu8BABj7WjcIlqe3bktTFiE1bQIHBuolLC8RgEiAaMm3MrUK4BhqnS9NZ0NkjWv0gbEmke9ipyQp3ZdtYS0cqsuWsLYnrulhZ/6qqyxBNm3J9ke3t4EZtQ49KLKolIkVZPv6gD3gkm+xTDnrUOPP8zNkjL118Unzb7u7vpTXAGNwJoGtIR3nFw+UyRlm8Qn+FmwBJ8lWs/gMQOI0wDBoDmYlYl/o6M9aEmBjTcFwdXt7S1/whGFOrQMr6hc67p1rQcwARVz9s/+5Ld12HrfgEQGD7+VeNcrDXjtDrfmMriY/01Z/69frw2vdy0ua/sigdeo+27x/Xm/wy7G6PzwkXpahmH2Oz6PIPdMU+gK5akDJaFl4UN1Ys2HBgJ4LqSv7Sj8UkLYbIFhATgaI9XJa4bClwKPN5vpsZ8lykcCXRSRgLH/bY4yyh87+vggo1vOtr6S9zGlpX/ZkLA3nsRDL17EprDExN4s6nn+7cKDNyifJ0tP2V+sXL9DrfnW6vaKPNfrgeuQR5BncC4jxRk6QstUm2y2vVge24eZ3DKbKvwMc+/jwuNpecdYZW9Lla1ao/7EBOf6OKulZQUA0edY8q9MDf8IemADZn/DkT9OnB6YHpgemB6YHpgemB/5/4IENgdwLYrgXBJfJIDNwNKA7eap1sh3U0jOXDCsN6szC8Jtg13AyoBQZF7RVsEwXPASojoJTZpLYZ9YSxfwTMYOcYQUduTmht0/Z/CNuJDgmCBUMsB6dUqVixE8xMJWRVz85UyzgDBkc6VN/tURuSCvLRVDN4HXsekKEMg2ah84QR18RBkr6BGOyDVLgq+RrvUUp+iABcXzmGKxSVX0zYmPPYktjRnA7gvnKPpNP8Sv79XXRaIs6WMpWwAgyrOITbQe4uH+8I9sFgEy74ZvD98e4+CJoSY1P9tgIzJt3aJw8dHBGUo9EbGm5XFvndCmr9dLOWhrVZt+i5Ewmm3DW2reEjr8jmUc2uzTMWLzGx7e3ZvLoN7OkSqP4HEXaDzQHHKs6HOJbfYb+yVDCL8pAKWf2E3uca/QV+CofFjiXdShjRi79oinW+yNFxrnlVCljLuSn3rGHe4Gk4mOLpbYt+xi5rXbpS+8vtpUspJScTMDQAS4nMpukPbJIl3quQVeLT8l1XWq/Z38VXbVHTflgk2+ybDAq6xBVyw6ll5071pd8RZsErw7xHfoOeeFz1r+e8fJvZd3Zb1Hn6A0fW8zDtN5niPlc+xthxqHZkQLOls7Uy5lv1LfIdRxfeRZjjzKol53Db65J6Sz2pV5+zpl81cOzbtYob6pkq6XP4M3pmt+yh9UTcqL64KtN6iBqFn+wzvo3sSwKKLa+5rixzga9uroCw11f89ZW0uVW93zKGUP2vEwPTA986oEJkH3qj1mbHpgemB6YHpgemB6YHpge+P49MELuCDKidXvlLdkOBnM5aD2BpfcGrRBUFtEATgiGk/2T4QbZIyAleCSmrFbu3YYogLARIPLcoYp3i4DvyBg17/2zJMg1IB/3uclXBcD2+2fJvUHrKPKxlitIRPjSZpHMILczy9LIV9Fm1JD9qS5NFyBhaYN2BVQqCnWhgU8BGBFoizrRlyv19hG35xLepWaCb+uW4nkmy82V4B53ITfTDFDh3fuPbAEbWVdRQSRKoIxwQ/uH/DCInuVfJ6V1M8Wm5yC6qsPwndlglvKfdsJ76JsO/JBMPXAAe8983capwfAJ+CFoZC/AaYAGtmXGVjNtbEfmC7N5omPZ3/oNVeAjr8taOLcrdpTohqDwWfAS2HAtO94SXrYhN9tzx/jnF+kc68ftxpbm0bTFYzwjWOOzUyBc0drvmL46LkBLM+BaPMuD9ql/tuvSp97tC6995lZspN/ryFg68+0+RXjvR76ta+vSsqSztG1efeulj6/ncamZtLb3tWnl7X3X7V/ySmWMr3uBN+7KXMZ5dmFOqstaEKhdAln2xZ6+OhSZMmiZbY/87YKU0nNdUFyvDXssjnWbJRsm478A/evb1QfXP8UMMm/1rTb5ESjzUP9sE6X9nuzNJzMjKQCKwcSvrwDcDgffYPkKPV/R9R2f86PLrYoN67mbZXpgemA1AbK5CKYHpgemB6YHpgemB6YHpgd+TA9s7h8+XpPhw8ecLUCuCgzZFmR4STYH5+nksH5qBzJ+jBY9N8tsi8SnaJ9A1UQtQAHHGLxzqeDTANUzigRrQpsL/RVou01OmQ24mP3UAW8NiBrntshFzlK29J2BZe5JlwqgL4CGdAIOjrUvwS6KmuW2A+RBEzAvDEFkFNIc7ym8oK5uVIexno1UGUrVXrLK5vTTLDiIphkXyFD/JOVFNxZgIm3ZCyW8u91B3bfkzajSg2+z1jggafXXf/Pb1dMTGWToxKhcK5AXKCv6AgboU54caEi2lelyVqNHZz1BMcC/kq2uYqmWAm6ScZQ6/g7zVJIBZMbY6urCVx08T8xsoA0ZZPEBayh0plQhWzkbtqgJkFl6DeTMLeYFOKXa4b0lq4n3BY4WaO0J3lBrR58Lrpz9po2st6xt/K9vVDnbBDPOVVMZTXA4y44OZUbarPuRb8Bj64ykSntnJ8GbeT5kf582jnnGf2ZFKU6WDKWQvWRmohX50tJ2Rqxt3CivbfGqDvunWtcC1GmLPyHWLtaWz0P0VwzFM8+yJvKM0gBNtfe8Fj/HVvvQx7eS4jMffYtAYumi5fId/ooT9Dw0AKENRGeOHdjzt1hXyeb0t4ISe70yMf1nqzrv0dkrTDPv0m9cNxTfamomIl3Dl3UvqJusMyeaInX7LvqbaWhBH3+vmL3Vyxskb/arD2SQ7XkD5eFwB0JW4/Zus3Rd87x5tFjWDjYfaL+7ewjvPI/8mERXWG95NSdqvAEofU3VH0C49QRQm2V6YHrgEw9MgOwTd8zK9MD0wPTA9MD0wPTA9MD0wPfsgYoWL0I4TXr3il1br4gStwaO2Sp44H2CRJzmXAgq2LYHIOpg2CsRYYJCg0HH1ZlkBQgY5NrPF399PlEJzVh7HG8YLyBF6XbvE3hnvLUqS+DIFuXmPKvR7/jwHOO8X/IcZKFpnW1rur522yVgH3zOnqsAXPoqfR012ovXCMAXVOqzzGAaXbmokzYu9bCj7W77bPM+9g/U4m95g2W2jJpRZuAf9xP4O15AjrkLf0Aqx4bXAELkZzm3n/XHn9IMMy72Fv0neg5fVFuYlQzaBR9Ln2rPQfUyHXpEFwi8us4EyA4H7SlfyFPdBU1ah/TBo1ZY6eN4C6PqatU2Xy2ofkNHm50DkQv5NX8IooOyWk4YhU3pII36F2u/Zdt9dW9dcG7jGViCP4j3mpclpK/sOPs7zOKi8BKgsi82c/X+uT7P6+phhlMX+4P7jYb2jQfhZx3oW0EhbLU0P8Gstj88pNN/lNZnO5Z78UQ3/5BXJd49y7BtqX/RaZsyy3Db/DRd6+ocR1fNwp9j9zKoE7LAmNRKP6+h6+IYi9Puh+/MVbY8astZT1gMWgHYjX5hq6zw5BOCbgFqHx/2qyvaTieyw9Ch9dPP++NuxX9R4D8cAJThx3vOHXvkg74YV2ePKR2vXQGkvUXWWypus6w0MxWrTzuO6izTA9MDEyCba2B6YHpgemB6YHpgemB6YHrgh/ZAQscSutnd3rx6s9lev+ENbuf/b1pBsrH9JXAVojDqtM3SAXOFyATWADMJQAVEoBIgOGS/UsgZOmLBcamEpBpj8NkfWoxeIyXB8hhn7GlwaoyrnAOBrP2Ky3lFyC+9S+eMRbRX6e3roFuNWn/vq/0CFNjmGD8ZP/xgu2CH9M23AST9U+0lEw7J4umMoOYZwIhKzlkySA9WFPgnWU2MjlyvbU/rEvlmwAkOaROZOgIqf/O730Z2GBiju9UREEEa9dBJ6laF8fpQcEG/U0mfjkTj0PvtUPqrXkAKFbnpvNo6m7o09gN0ZhC3lALX3FIJT19V6FldzJRv14x8D+LP3DCeBumvsOfaNwA+1XoInwECVsZeywJMi25DxXGuVc+V4wRUfKNjtgCrH4BMzr2jTy6CZHmjJTqFmPWqv3pu5RH/SEzpufAaMEqZMeSSdZc5QRQYScaGFw4zA7Pm4sJL3uHrfAfwKXA6rlTeYp1J2/LP+o3nwjexdrHPzDGLb5a1fgZk0TUy9Yk2CH9jQzI5RxZhBh55C2rmpehJqKo6+aWuWSxBt9EHn15HjpWvRVvb3uKVRuaj+sTy7E8fsvJM6UvJ0Ln55Oy58Zyf1nVuG++jgB5fKdvHB93Di/k7Z9PhRJ8o+fsCC/thq1NrrStn6Ji3flI/Ypl6XPtMoeDNlVezZ5/MBMsSSVaePuXzCDh2w8H9ZtWavVm+9uFDv+EHVuk18/BTzP0aEddoSkpaipM/VtZomZfpgemBucVyroHpgemB6YHpgemB6YHpgemBH9QDzwOz3dXN7ZfEoF8SMF4lcDZ6TUxc8ZuBpMXsHgPOOpiaAJO/gF4EnvYFkLC/A3TGJdDtrVDUHe/HMF4yQS+vtrWcBpCUuWy333oC49xXkCudfQV2WHvWvgjam59XA9ozT/R3+1S3q7f3Xfpe+vJG9dhuS7WXvbWF82Kr4If8WpaAhaX5hMdoE6yy3TYD7x4Xevqil5XMYul3JKj/5ttvwTmsi0CULMkwkskZdhTjAAeti7CAJXIGWetjmz7qunS592YU+dAog+A6R1DPtAmWUYLhCOCgm7MOrBGeWu+bL+UXcMQXDACYXV/v2NILePNYcyOvpR7Sd6l7eaKjf/RJ71/xtVUApzK+oo9fybDTGdxCL8vSrOvFxzUdfqHx/oBuV4AhjXFc/NF0uCH2aF+3+fZIbXR861VyF2t+2NXt6qbvMy+Rf1mv3bak9X5ZnHbXYQBlfHD04ex1CCgmMLYjEys8xlwJAlkayG6eysMc5hLAKLBarYmAZDG45sixvV68bz2X97gA8HDM09DZMRblRda4z88Gegp1HRw42s2MuwKBfAKgUoe8/AIFBaIF5OWzxbb2XxArf2/yfJRe9rWuAokCp5lv6ZBn5ix4W0Cy4+lq9cD5fk/0udWz/eL1CXn+XHoG2T1vsjxsr0lw45cIkE3QjBdn3D4dd7+E9pcwvmVFfjtmCu56dZbpgemBpQfO/5Vu2TjvpwemB6YHpgemB6YHpgemB6YHvkcPXFAGEpnuP354/eqL/WuAg11nnRDQGScngPMAa4PBxMlErcG0qBNWJvD3mn7O5bEcx94u25aAQNfNrrmEhgbLBNwEnpzWk/El6wLyZHsUvPhHgZ7gNrxgYuaY8bVv47N0sN1gSdoS9EIztnKGkK9LAF9AwnnLHQYKmKikYF0iWcGGUuCZ7tDwJ7ngVm7KjOgb+81wgaO8Su/SQG85IueUwT92EqiLZajbGiDBLDkBghTGB5wEbBnOWPGWvNX7h4fVN9+8i6+jAnRJYSJyN5NF2aGnU04mc1l4TWndVMWW6Gf14pvSMSRoItinTSp+FP2KavI3s892tB12lo7OI6OdM8fFrlpYnm3ndra1BlsABN9+8VXOvHt0UikCSwyubDGaAmaJZdJ/hfzl+qoMIHUoOwqIUbewCq23zoFK+RbGyii7ADOxrcizlqzXmxvLJ3aVzLEG6e/1arv3Z/6I+cSPJZZGddQq/YAe6sJYaZt/87Se+fM6eHuNDmM+AkjDEsZgYOoF7wA3PhuMJiMsBblmQ50G8PqUjClW73acTRb9Lrq0PSJAuQci8lqAX4FIxRjJbEm0z+I1n7FWvN/va30UoD70p915ZEToc6Zbr0l1RJ8s9fiFCsUD89eH9eppXbq4crYBgLHTPngK1fo75lrTe5kP2uJ0v+lTe5uOA3hzzbhGLfpPuTeAXOXzXebq+OhOZXdI+qvjK0jMiKzD+u/YXulO1PXVGs2YUvQf83rLb9KveInlr1CuDteLlChUAqs+v6cHpgfwwATI5jKYHpgemB6YHpgemB6YHpge+CE9UFFsJBo0bsApdr5h7RWBXN5iaaBO9gN4VYFOkhp4NviUyNXA3kCUaLIzugz2i7bpU824BK7wrYDTdsP+Ap/sS4uBKbddTyNfCW0Zm+1W1Cvgrau6FjD1aXuPlfa8e2xYLn8/2SYXwgJIwmvoEh2MlCnyyJjULnJG9axP1/VTy1iOs7/5Nk/blvbgkspkQeaZBjW8V5uMz1WvVPEcpPcf7+mnLS9CGP4cAb88hQQiR/u0i6tgl6W3yMV0QaMhu+WfBLCGX0LveMuizWromQ+LwJaHuQf+gFz8oUv0oKL/pa6MOqGO4+rLN6/O62yP/stxzo+rRvHew5VPlfaLNe+V0fNgW3TzKjjCsm7VowusBB6XW2Ed03wiD02VGDkCgIIhg0lfHWNxy14XdShdS+dkdLX/pIXH8tO+sS06j/5eq7Y1TfcLuFW7vqE/c3hZg7apg1tx8wzjVNdMnzfWh5UJNDVt66QdrYs/B94LKnkVdpPezCugJGdGct/ieLap+4uvW2tr7Kdzp2c/LfIPO/x8ZGtn0HrtZOttz4MkaUcHyxagz3Fr5Mdf2Omv1HI+pJNGfbwWmF84lZlgFgF7i79rgmS+tVSbHhZbT+W/5j8IeP7ZE2AY/7iyRXN/tX46Pq1vb29PtK9vtsdrfP4Ttth+BeMrBrTpPhGLpyIi59f0wJ+8ByZA9ie/BKYDpgemB6YHpgemB6YHpgd+cA/wgjmzLAg1t7sNYNgtAdwtQfQ2AT2Q0xXR8og7CSQLKDNDx0LImYA7GThpMIDlxoDUgJn+vFWOgDbd6SxAJFsxzRqize4Eztwne4pg035LAljiXmGhAiNoNGOJkkA8vC/xZcuVr2ckWWxbXocakW27oEHRmClCw9h6Z4aMDd3vYeZ21zd2YF+NE9xALYEm0+0C2kjXfEsHbUhQTmzsldaqI0M+8s620iiBffghZfT3eUancZ7byUy7Yfpmd7169+Hd6rsPH+BZGS9AnkO/YpPofeg2WmKf96VP6RSb6vbT8edBRR9oEzsaYEu22qAxc6Z0KwCmTNKfEOCnDWDH0XUn2NHZOwJw9jPRb7/4kp2WbGU7n9llh+fskzE2AByBC1YYusOHkjXrXAIM0egEMBesL+sM74Vcc1Y2mG20FXiJsiUjzMZXz31Va771VbYED5rM3QDcch/wp3SS1mfMEpf2XNrOp+c4ciTw44U+n5/cx0e1Vmx35aMJYF5lfGmbQI3LJbKGGeoivdsN7duwLXQ81/gcLmYpYr8rL9uBeUOH9CcysyyHzXg+hb3SBD3X9WOBYQ04ZQwMNz7Pe+yCt217Pl61LQU7Uk8mZ61tuqOL7fkhgLAzJdNG/XytIamr/3IezW5VTrZHAvo5RkDN7EQupT/K9xpRnzUd/qZkPerR4bf8rkjgOsU3+lRf37Dt18w1eerv2sapY8zYgzcftlKuPpJFxon9q83NDQf270++QOTAjwljXjw+3b9kQF6CogjncpbpgemBP/TABMj+0CezZXpgemB6YHpgemB6YHpgeuB79kCwCQCVX/6dv7f94ou3twTKt6fjntwXEY4Ep+AKBeCcg/kR8P8x1c4BrQAGgapB5eCVoNZANoEqQEfTVuBawI5tCX4Nmimh8ZZPztca+tiXDI5B3wFzX+33vvmNMN3mtHV715s28kQdAhyU7d3XtF6NqItW+7AFATSV7ragb/WPtjLHkUUz6s07QJNiBS5ENNymuPCB903b7frSe4GBO7LHDoAc2cKos0YJsKbPFm3pkjdywld5z4CcbJGsqUMnbS3ATx1iaOytdvmpuqX4AaICyIiphp5zxdbbGztT1z48lnv7N+gv/+OB/WssytsX1+ED5AFHwAhlUtpe780aiiz6vPp5XsJ76F1jlMoftro9bjku21jxZ/QdjDIP3J/pkCE45jZcs4kEYTzbTTedD8HnXh6q7LjoAL0NpWPZsuQ9xJ0vGQdAU/Q0izpRAgChv6W3xpasCAuoo1zbBEqVYUbYdnsFuFiA2mB1BqZ9hor+jZcjjwAAIABJREFUMh/yd9tjyde+8pUAmYlxGcM456Pta3sCLKvfmA+v0jUAxr5D6q2jksa8DQCt9etxzTc8JE+pdV8ySjeBVmkB9SO73o65P28Fdc4DQA8O4rEWebT9jsdzaUedFDNWlX18ghe83c7senSMH33BV/i4qn3L7w4UN4AZh5MB0fH+hDVqcTAZB/TzfKs8DogCQ0rJmt/TA9MD5YEJkM2VMD0wPTA9MD0wPTA9MD0wPfCDeoDAkFh0t/oP/tE/Xv2X/+S/2qyvdjeP+/1N3sRm6EeEaQDYW6UMsA0m12RKJKgckaznNxnvpS/BpnUj4BE8V2yfDKuMg6dXCGJvj7Pe7XW1G7AoOSXIhKUZL5ZktBCIEmkGmFDPHpMQF/b99j/usGZf2S/I5dzuhMCOkb8Xx/pmvvCIPRW3GmxH3pCZMWaLCB6gz6WY0VM6oGkCZ6XIL2er6R8zTQp3HO3YER3qKpARMEDdgyA0WFO6SOunM6ba3pw9RTT/+2/frTwDSRcJOIUePRmggIBCORPJukXZ3Yc8uFez303DHAcckM8oZTd2edjSYpzAnnOeMsaXfSXHe+dEsZb0aSfrKvOqjqjmmWtff/0TmuuNgP8ve+8Sa1uWpWftc/Z53ke8MjLyEVUVrkyXCzBINArLJVNSFQ0kcBMJgSwettwAuYEQHTo0EBISWLIEPQuJh0BCRiCDkOiAkGUJF5TqYSNwCfJBVhURGRnvuDfuvee5D9/3jzn2XvfEjbgRWZVJo+a8ufZaa84xxxjzn3OdzPHnWHOln3MoTYMf7UnjUNp0ucblWZ99XVJvxCdfusRu2awMyCJQeq52/V0v3LHGRMROrrLxD5zdK65t2eIG8ReumYyJZwRSr7+i2L51Rp39PPSjdciThLhhqWVdZR3WK5ni4roUN8sGonGfTfQlQX2hMQQxTWbTud+Ya99XWtXvypWsCkHNMDIq9cByhWjDZ+257tQTXeKPbkttes8ZrRk99aA6xub6r3GIQcaXXuA9/i7s5zXfGpu+iVvKDdvcD3JqdMl83YwMNj0tnGqh1PV4NjKKLLvuGv/NNPRLrpkDMg8dn8NwrdzA6ElqymVmaFynjPWQNUFFZhDs9iHExOVy/K2pV8eLnFxLMjK+wqjOyu6Dd+3zRn4t9i/PL2/cpJ8va+6xSd7+3sEhU7Z3fnl2fiGg8XPrRV3M34nARGCHwCTIdljMq4nARGAiMBGYCEwEJgITgZ84AoR5khkEzH/pL/8rqxdeefXgw48eHN/ckOVAAMnrbbwpWAQNAeSIKA2aiSqJMg0Qm1CpYLEctt2j+lZdZO23KNYZrHab8nTcSkRPwluD4TLfWUT6B6OylW0dXeG9xcDV0v50xlGRNOVn+xDBxY+kID3jn/qSJUKNJEOyqXTXa0q/ambYW7bLvm36oA19yOtsnNs/67pkvNzG1iAil3goVwTGTrd19pOogNtcPfrkyeriHPKHOVXPBtIgRQfaW2RvLiU3nPuhq90QL+tDM9hz56v6bvtbsnYZ60RiI/3tW2Nx3zL3gtKE+GdOuFdfMsZKMPchpHylEmLs/r27W8wVCY7RAdHR9gaW7Zvr0evI93hzB3bIFtVZFZGDAOEzg1Q0AF46hsZFjJSpeW3d4qAPvmqnX5KekkxmDllqLpEZvrhWC5dd+1JX4934evZrk+rutR/FPA95TriRAHI1et9r0/Xi7ImjOvMPHyTY1HXIWLXrq5WOy6cjY+WjFT0eqqJPH5Rtn1zj6WtX1Kd+4BRz6hrjtS0EXAimWhvq1QfLAZlc7bN2lbet9NfZOppSnq4vHTZY3/29bx3Oqa8/Qk5Ry9j5pz7lPVvs532XItWr3fq0lWj5jWhhBJ7MN2lg3EOEIaMZtGETEh735I3JBr25uLi8OT4+3D89PHUvxydH946+/+jRJ9/F5idtl7MDGpYWtfNyIvDHHIFJkP0xXwBz+BOBicBEYCIwEZgITAR++gjwP0F57e2dd95Zvfb6z7Ivzt4RAeShfvC1NSLKCsh7j6lk4QwnE+yOANkg3nuDRItheoLoIZu8DoNRYvoEqOg1QN6XoDMQNnA1swoRA9PKgBm2DWwJH3cUnUq1Qx/sGFnWq4mhBp4KhNWlPQPtERfbGQ6k+q8hLozhfX3M4NdxuE9VE2jeu+eVr9MZ8DvG2NMnx7NQmuA8FEzZ1E68Q2xL7FlJScYXfTtYr9odgbD21TjxGARBtxfpQD90xj4Nhdf+6oLgPK/Q+cU96j1o5GLE34yBV2epg7wYxI4iFZ/XlSROvVZXVFL2UnOsAT8aI5gvDqLbZCTHEFS8gSAMJJBFTlHGp85UDlyG79a5B1SX2OXGzDf1HEmikA2HeMboODv7zj6ZLxF2Dgd546jVW//sqCRl53rdW6V98ZGfGISiwO7qh2jWqGNlfYz1a7fGPTrwlQWd9RE/1a1m1kva24+h0jrtSMY5bseii51BBe0yfFMHB3ZV0dmMrVfCUSLogEwt667HfKi7CLQapx8dcP88l2e+/ug6lxhkQE1UhQMXS/uSoRYfWYNLPLx2xjpDzeFYd1tmuU6V8fnNGMdDLH6SixLd9g3BBAbuI6Y/63XtnTfE80xKpgZLkKizM4dilPu8Wuc/r82yi4wTBi7MQvDQVhXqqNcvi89/9mDj3r8Nrvd8Jbaai4unrdYcG/Wz959fXc099Ye8Snwj6StuzIU86Xr/AI4TSpzpRXR1cHzw4dHx/q9fnD/6O1j5YKj2JIt9a4UsWuflROCPKQKTIPtjOvFz2BOBicBEYCIwEZgITAT+f0KAMM5CRgQbvBNorwlOD27Wh0SnBNTJrqkAmJuSNLKldKCZkHQE+wakFZwOUgA565bBs0GppFuCYkkBM2uGzvQfAXPr9z2kBLHU60PL7vZ6qrrWl9f0hn9L27Z71Ct5RebZ7mhil6C6bbYNmqoNP2vUNe5qlyYQkzE+hW+V6IvbA2baywe1lT92aXu7tp1cj7N9MyAvDAexIIaQae4v5X5TP/rRu9hgXJiQaFB3ps4KLzwP262z7Jc/yVZCZ4amc+nsyXadLX93I/r0Pe9Hlt3Yoh1hX30L4SApQTtMF0RCvQaoGb2yxBdIGXYzX90/PQkhxU7vEBTYV0jfXEOjbLEbY9Jk1eUifj8lOxx3PGLZxfvWVfVlo7B0XRfeEnQSZRJTdtfedk5Q1hllrVedfVgnhmVnZ8/7nqvOOLOu58d+vvKcjeEhurSrzZYJEcZzpA5Xqv1C/qhjQNWEln32wc92ny1fjba/9c6TffvQ7j7vItt2FeKsiDzrHUf717aqvnDNGrW/ZBP9GXXkvbZfMtoGdq0HjfHF/b3Ub2n5bstrlIy92yWuu7+YeO1hvxz6mbXhsqm/SzVf+lY2Wt67+nujnp7/4Qj+By9kfLXV9XxE09XVecjzDa9v32z0m3lwHIfHwYyxJAtX3Xub6+8dHxz8+uNPPv673J7h34Hucu3Lpm2Iy1kmAhMBEZgE2VwHE4GJwERgIjARmAhMBCYCPyUEmhwgeYHMI+PB6w0hI589NNB2Lx1zKvgfqMRxBJsSVItikJlCmyUkFudNbTptTQJUFZtcQ8hagWteeSLANOAcQTqXWwIiGWrRWZkqBpw0aiL9UVp6Rn/JNsWppd5rglvuoWBGQFx+FtFh4BtN8c1xSdp47iDZczJIELM+eybZZwx3O24sRHb0zwjVg6ieN9FhJok21eV4k0mnTDnCVV379Uv7iPOyzZENjiP1zkuRfGXfzJT9Q7Ktjngrlr7f+c53Vld+QW9k1ESXmS3iI4xxkDuU6hNORa99M54YU3D4qIwH/ganXDqoktG/skEH5bIuVOKka6zshDARQ2Sih3HIC4QsUydABSPWzyFr5ISvBb7yMl+xxD/eE60PDyQPiG7YsN65uIaYyDiojv/6FT84YQNUS3adAW9lkylXE5O6+MR95oD+1aSv5X+tRow4Xn3KOJBnoSnTxdcQXa5mITpzrrvgY8+FoNdtM37naWMM7N3uuLRPD9afuDhkwHOuuNnA1PBd2awVq6OH+VbGa59fnwAxktRpferU1j7ZTw7BdX495tHnN48mPbP+6aes4/B8NHR7nT3QyJLqMWSO6Oc5+nXqVlG2/bMpzz+z05lmrcO2roscurpN3SEDaWi/4o8AiRWyvlrqWJJt5rOCjfZTWduSqcofJXGsUv3NXgM85sC/fYxHPaWZC8dkZw7rsLkXchHykDp1WyTOqucGF3jpFhIMv64Pj9Zv3r17/Nt3jg5/9/LsyZmy9FEpMzHLRGAi8CwEJkH2LFRm3URgIjARmAhMBCYCE4GJwE8WAUiJ09O78hC8Yule3xAPZo4k4K2gdw0T0Fku5YxBoQHkCPRHIGqbwaI6DGwNJKvOGNMAU8LAmLD6RQl3LZsgNsGnG5AjblA6SvxCtzqvff2QUtdSeUVh4G3qW492LPpaZy+KtGgZdfRX6lqmCRQJq/i21bPzR1l9Sn8zSDRS5upaAYrttlV7XTcJ0MF/y+jHsk/pls2ocW/bIlU/yuiH5fGjJ+WD9rhvvWlc/IRH6ntki3gbzo/6Z/aVWcFel4yJ/mXMOSk/0lch5DNT+LfmNTRog8Jz6NiEzEFuEBASThuypQ6PD1bHx8eYAlebkY+ZwKO9XATT9rPxdQ1IhFiW6ydzgB7JmSJTGQf33d9z+qB7WWe/bouAPxKzaDpkfVxKksEzO6e+4prmoVf9ltiOz0V+SUhm7dCWjw4AUq+ldOAnNhfjVLWkjPX27+K96/V2KTnXnbK1/iSBMh76Zw2YzUeRTGxyNmupAbQN/TsMtH8cnbHrVEjGDr3KWdy/L38vqF/2F3vvLZ77edX9xqj8jUhk+lmx3YC5nxnP+mq9RLRF1daHEuZ6mIqMslt7LkrbB2ztY/400dQ2nGOLNlz6IeCitP7G2c/RmDlLa/+N3EjgkSWXv6Vk/n0MHr/JW8f/61u/990fvv2D76tQnXoxPOdqlonAROApBCZB9hQc82YiMBGYCEwEJgITgYnAROCngwCBI5u2E0DCjG3YOIcwkqyyEVUmgLMuwaCBnUEhh9RHAlGDa7MvPFNvFpj7dnlNGJkhcJlIMNkdBskjsEVFgtEO8I0YJeY6U8Q9ygxBsRp3sBB9vqLlq0wGmhb7dTGYNbCNj+iqopx9+9wEnnpp0Vf74Zcl19SZEXc7e862/lqluSb295VUL7RQ424dfW5CpLFLp8ItBmN0O05pi/hPDG2wzY1SRuL4VHacLmXEyuPR2fnq/IrssWCODG0hLsAgWU/q8RAt1CXYD+D6tPNTM+FUUukdhYnLuLZZN/jlHJr5NTBz/ouL4exrkqwJpEb/wpcW7sVMnPEdIkyCKEX3+PqfPvqaneO7vKzXBvMVRoQkeK4Yo19mRAANrEKY3f5aovgMi8me0lzhpF0KeLp+re85troz/pTKOK1zfPjmvWV5dn2ZfSjuynlcs1b06zpM1tDf3uCu5Iya1OM4fKbSN8SXeBQOsZ952vko/bt8TVJ/XHu9znt+rG+iyzNbYCGDVVRrK+34qO080ww4z6644VeeNs5i42FHybhaJsiwmX90QIBF3nGhK/OupYGr3h2RBdgYq0r7dR8V9N9hmpl0rSOj3m3BdvwINPjhfIC5dezxhZUah0Rl/KDe1y79YqZ62obyfQRz98ijKBP9wyDMVq62vnKHSeYWecbqOf+Qs59ya20xn2sI3bP4syIXl9xTCLLj0+PVnTt3HpBY9ncfP/jwd/7b/+w/+vjqvTfR6rZjLFxc4JhlIjAReAYCkyB7BiizaiIwEZgITAQmAhOBicBE4CeNwCbZOjebPTLIfKtyF0wbBCZgHYGvQbcETQLVEZR2kCn5caAc/dPnttuSXWTAWNTrYen+2zNBp4FnCJch223aqFcMhw2C09ajrmddW9f+9FnZzypt67asY7ZYb1QbOV6J69LyJWdw7lGtnaFVPbtH+dv9rNXX+Mv4l2NpmR5L9sKK/rLjq12Xn1yvHj16hBL8hASJLnwWy+zNVk5jpbxo/aW7MAohJPbPKC2fph5Yn1veOb1dlzZf2y2SMK/9SXBBKuR1wCEv4SPxeXV5teKVtJBPhWGN0f6ST13nvk8swdxnPaKn8enXZHUndfjgudt16TamtmXdjbboVJBim8U+fS2pJtl2TGacXw61TZyXOuyjvON04/lkno25dazK1n5mklbiUzaWdsrebg2rM68GQ9bY1mO3j4dl23/c0zv1LX8AyYRDIScl+ZrILH6oyDgeQPQMQizPnXR33ausfB82mYjYliTFJ69t97rv+7z0N4SvpBf/JEWvN2QPugWii4TiHmmoYDnXK6Pq1YP210fSuqVO7XQRd/3w6OJTLAnfPnruPn3d9xvmyC9+qrHr+hxy1C+ukhl7hM/XgHd+fr66uLgwgy7/3wB79q/2ri/eg8z73Xfe/P3vXv3oTdjhaz6CAlDFku2cbQfneSIwEQgCkyCbC2EiMBGYCEwEJgITgYnAROCnjECRPmYeEYMaSrJR/5V7qFsINUc2l4E/YSJ8VAJLg0S5ro7uPBtcJpqtrtwbIC/k026jwW8F0dGzCFC9N9jN1xMrRo5e63aFvjIj6I4swXRlsKBZv7RjLkzORajot8UxtI0KhivQt678cgjoGLL2OxzBNRpjJ8E4MpJJpXY4qgFqDMZD/CAvwRB9EdF246GslWJaWS/5YEH6GPBLuFSWjiPvTKayp89FGJhFp9w+XyR85523Vk+enNMIhdB2GPG2aFwcmcsbyCnyXGji2vrowV98z336UzuGZm7Rrr4q9VeCI/XBmlv8z4b6OoDezmbSh8Kbevpt/HqlWYsQC1EDn+BZ0otlszo5Ocm+apvzh8lSKx9px38+DcgrmCfIOU+1Xli3DoH/8ENxL6+ch/8SLuqVjJKIC/LJYhNLfRBHxoj+kCneo8BrbddaisrSS12TLp5DMjkuPaCt5pb+AJh9zSSzxgb/eb3zkPkDO/uSbBSf/HKkGZld9MkvejrmfebYrChTtNRvP18+DV1FnVmb19c8w4zFtoxTN3w2kKd7iq45J/VVUjgyGRy8NlOz+nHPf2IvwuWPZN7NyJBTn+vCKfdYQ85qyrJmXDX+uo8yLrPvF4rtp7yl5BwjlSl8LdYvW1Iytyh3PJHDP58p669cN6MLQ49t91WzvXUeLDL0SjWCjluHx7iUDbbgJadcvhZeeBVditIxbc5te0orY1HWjEck0OGfTD8i8OjBw332GdvbP2atXh865N8/2tv7g3f/4AewxBeYuRYwxNUbw5xnmQhMBG4jMAmy24jM+4nARGAiMBGYCEwEJgITgZ80AgkB3aHbOA9jbixNoNp7ju3fGHj62pKBZRMFnj16zywjZYNgg36D9QShep4MENVaRdhpG8WAsoNTz12s76L+lmu7NxAo2lyvjxDTY4N9e9QwWi41Fd1Wts1gCCRAuiirTxVUV237ZLDsta9ztX+xQx/7eaS+zA6VdSNeCZgTsKMJ2dsl/fEZTcGqbXi2b9sIMYbafo3RWSp/nx7vev9w9d77H5bPXMs2RQ71GbJhuiW+m8lEf+zcENBbh3CdEWnMI++PGI2bHssWs0U/RST22Kk88xL9tstmYCNjYXpDRClM3Ub7YuwrmeIBU7G5OGeTfl6xTLfCWnGL9vWvSK5aQ9XCr2uBk9ljIe9sQD4+44Y+JyMqzK7XjrnWW4/LLsvifNxu815dhW+TXBJMvjq5fW7ST5meU/V2v65zLBJkZp7Zd0mQlZ1aS20T09EhqZrXVFlj7ANPZcm1DSoiJ9b21V6XrK9BDm6XhZZVLjauSnzK683U7fxQJq1RFXml41PJdZ0C1a9WjkSfpe01rsp4tH/6ZskcM8ZlSRv+HRxCRuGmWPpcpC8+WJSJbtcS88tv6rVR+4R56xgLl7YXofFj/yVBZl/xtmTOh5zL55CswEv0SYztHR3xt/Jmjwyy7Pd/9/j47PLi/Pv7Bzf/x9nD995987u/i1ls5x1c6eBZJgITgc9DYBJkn4fObJsITAQmAhOBicBEYCIwEfgJIEDAJolFpsl6beR5lQi1szHMdsmG4MokaDbwNGAsV7y2GCzS4E/aKnusw9NNAloTm4gwE2TWVyXNNqlX02jZltZpRQfOHZjalmwdglIzahLMGnUPIsA+kZVdodRrayMLZRGT2sXX1AiTo6MDaz9G0MXNx41ns4+XQbXEy/Df166kE/cr0y4BdGURFcGl/nzRzv74bHzdfXPWv3Ix7V4mw2jgqXLHJtnoxvbOh2lAZtvYv/d4k7hcHxwlQ+j9Dz9aXbDBPQwCyrQLoTEIh417yo0S32hP1hTt6qu5K4HGPHfdhojFfcvqok7acXCO0WNjZloICPxkTcUxRdUz5iTkln45aOq8vL5iPs3GkTCjvHj/Hq9b0k0mxAM8XCuxpSqOPV+3bKJHs9iQHIsMc+e48KiIEaolVlUV6LU9illA+m6puarxjObo6TbP0TvGWzKQaDiUQ5v6EUJKnYWLcq3bdWLxGZA42lvz+mXv7TX8yDjoTmJd1oHyWaPtK/rjMzqueSXVjMsb9CTrjOsiorGNL+mLHzXPjk2vqh6J6Ekd9dlwnxufC+kl51JdG/3jHFIxGp0RZHwOkAsRF7zVWGO1PjclUbiVWWczWrJXmAuAuTR7zOzAjMu1o+88j+rLgyiuqsQPk9BCzrvG9Q83jkLqX8aXKyaav2esk8oqc45rPUiMhf7KuGoMMbO6pE8w0p6GRsm+Y3HHccYbWgo3feZblasL+vKMCsbqkP93wQy2w4O9j8kg/K3VxePf+q3/+X/46OrN76HX59g/pkpG3ItZJgITgWcg4J/1WSYCE4GJwERgIjARmAhMBCYCP3UEDNrZCP2AADDRu4FgB4MGjUVEGaDWdTvYAWXLWm9dHxVPEpAmvt7p7P7LswRA61vWe22bx7LoU4ijUbns29f65XXzOor22Nrntrut72yaIdt9PFviB8RM75PU/ZpYir0RSHt9u77lYR1Kn79ct8+p5Kf9C1lJXO69Mq1fP3pe5BM++OCD+LbOa2pUDELKL0XuyShIXtX07nwKkbOz1bY9t30udtXYX7Ztx7KTqCvl4AFCElqDg9GHD/v41+Pw7PhCTNIle2Pxuu8dNjd3bI6x/fDsJvjLOlW3D2Jg0UP1dmn8W+52/5Zb2um65Xnpc1/bR30+P0WW1Kb91ivTOpVZFmG3Td+WMl57VF/mmjnsOvu3npaxv7qUh1tSIjqr/mkCRmK0dXluv732FcrUDUar5ZTxWhKoSa2Wiy+OMVadm906UaZLj0UISi9/D4begoWsMO8XeDV5JJkaAp+2Z5VkutFX/yS+nAd1OxdLH3INlvrSpa7Bf1tV86Vsy7ECt9fLfjUm9k0bhLr2qIM3v7465DXTu6d8sfX6/OHd0/XvnH/83m+//92//+Hq+gzF1wLjTD09Oa18nicCE4EtAjODbAvFvJgITAQmAhOBicBEYCIwEfgpIGAOCyFjZWEQWLJVTjEoTTzVpuPEdfxbG8SOzIlsh0QgaSpENoAfAX+CaEJAoz8DzaRKGBJKBnFWT4LVhNWVseG9eSK+FuernctSsqXLoJTQl8CTfuqi3wGvE1Z8W3UwCqXfTJvojNktEdH69MdAWt872I1dSB3rpAOUdY8vI+gO3hPV4ke+lAczYaSr/ehakB0BgIZlvdfbr19GkaRJea9t283Ys+iTJZl6kiRe88/MKdv8F2JJQgDIlP7w448LcxkTXrsLpVEZK9HreMQs2ryOnJrpr1nqOm5XtskbCYTyRkGB5z9ihL+Wxi8+q2jU26aOEHMSDbGHvCQZTpvt1KXXW87Yvnd8Cr/X5GKddU+/Gie7HwwCqbLhxlho8ErZwgC0ZM/QJ+GUNV2i8R2HkStfxCfF9cN1srwYj69+ZnxutL8otQKwM/zSN0kaN4HP2ljgYf/ynfWDfLBBl/UeGXuInszQtj5fGx0ZcQwinkYClxFnHiprkw6rmwszscDajDb9p13dXktCeg0AdJJ89Ll3MGjj2r8EeS2R89o1L1a0WTLT1tHBZ6LIMFqbsCz4mpNFt3Nf8prEi/IDO5b4piv6WAJ1HtcI0MNR2i7+uu1guaBNr8TZwhObbLA95tjubvFl1qt49ldcHYFt4p8Mv2gYPoEFvWI/8+Bc204H74OhazcF2/HZ8THHrBNxNGONP50sHzrwoYEjknEhyh68/tWXvvt3/t7/8v8yMTh8cxxBcv4czVA4TxOBicBnIFD/DfMZjbN6IjARmAhMBCYCE4GJwERgIvBHjIBBmpG/webh3ubmDgEh7+dVIDnORqUGf96mGDSG0OJsMejsYpvF9ucVZROwGvByNHmwJA68Vs52S+vP63JXFcAq0+3KVABbbd2n7XhvaVteK7/sb9uufkcwWLe1D3PV156X1/rTY3iWb61n2cc6S/vhOWH7GLd6lE87hMFyPGV/tXrw4BPaJT2YK8kNY3x+WufSnkH/U/bGmFvvU7LYtbT91nf7nNcCF2shnaSJ0l+6aFeCj+NBtXrarplMkAiru/dO4XDKbttZvgopcVXjbhINPci3j22px+F9XddaUWev6dbfGC91LNt2OkrXVjcEyyF4d/ZSj6Vs7Nat9fbx2Wi9kobalcyxrc++apiCXkkeS4i3+F06W0caFz/sg5VsstYbubGOpAL1w83vu7/n7VjQ0/63yibDzN5Ttv33umW7//K+9Vun74VPjcO6lu3rvo9ddEvWWbIRvudQjqnKjzaVKTkJv53v1kXvAms7qVJ87NtryHpxz+vMzIVliwlzO9xInV7U2q1MvX7W4jsMHqTu3vHRAV82Xd+8dPfkB1cP3n3r+//7b7Gmz+jKK8Ih42Ji/kwEJgLPQeDp/zviOcKzeSIwEZgITAT1l9hcAAAgAElEQVQmAhOBicBEYCLwh0WAcI9I0t+rU15TOt273jtM8Egwyo5GRI5FKJgxZUAp71XBJW0E7sSxFIJUAmD3i9qnLgGkdQShpp7YzQDSfhZfizKxxiwkcj1KH/WRoZ9n3TKgjkmMdN+yPbJtcAZp5CWTRiCba4PmIvSyZ5ZOYrp0DP36MfRWfY1Tak//48OQkZ5o+4UD/huY559CklcG1j3GIkDs0zaS/SJ424C72ja8cWUGivlhXSQCrkcmnJC1HqGu1zoHjvivfjfod+uujx6QQUYGXu3NVASEWXnJ9lKPBiQAoog709G8VY9ZM7SBQu7bF4k2+0kSKGeJPz2fNAQbiS2dLRHmGCyUtzM+pFlyQNZOoy4MfWefKHOttC3BlbVD3/v379PMPQqami07ZT+21EFxPdG1SmzWTc9jxocS9yvbZ5yKBAYHRQnxhs3CcqxHF17aal0wS9xVXRrSNtYACl0va7886qbtOHPlWMFDSJIGeOB8u7rKjmNzXhxTPS9FlGnWMcdnDUHmqNujsGF+9KMHbD1i/Xpj7NF/3w81qAk558H+tmnX1wJ5nZp7xzPGR33Nr3XK1Too7Q7CZ7Hkm6jLfAxZ27z30NayLOXKhnMBPFlbhUH5ViSj4wyxyzjtG6t7ZvSp1Y6ewNuxJ4NLTOu5dZ5u2BjQ9eT+aNoT82S52g19vg5JK+vGvxs1D2rWrkSZhdr09RERo2txHOMq2Krda/Zo2xyy4dg1Jz8ucefw8NHV3uHff+n49Df+u//8P3nv/K3voND1cIE5WP2sDfXOMhGYCHweAk//Jfk8ydk2EZgITAQmAhOBicBEYCIwEfjxEUioSXfDP4K2BLZ3CR7vcZ8MMgNegkt4jvqfqAaWfSzNkjDBLYEmwWWCeAJ6SxvIDT8JeiUnJMfQZdkGy2Ur9eqw3qPt9XX3kQCyrfu3XJTyo46u677at3RbbvhpHX3+LL3L9talDuVzT8Be5emRtx+jMScha7+sKGxqTF63re4DIrm0vg7YHuJ4SQEzgbhaXUCQnZ9dcEUdpFMThAnGlaCvY+ci163bc48h7eN+2f68662/ZjqNeVEnA6sVliXG/WLOWmdnTLl5uURVPggB0XTv3p0WYZHWfIZU29bWRews6hojq3que3zWee1hW/vd52V7Xz+rrXUo00SVG9m7f5oElASSX1rURh+tr9ZKrX+JqkzJeCbUG5XgplxkU1N+ty/KeV33tTbc7B5GaNTzKi9Ej5lSFuXVVfr3Q465PkpH048lp7z1ypa8NYVl2av7ZXvL3SbOrLePGLSOZ42p58Jz9ynfyg/7to3dOOq56Wej27ufupwPzx7tm+1iYz+vW7d6PZZ1aRw/0eO1pNtYzz5ro7DN3/WV/wfBnZPj1b2T44++8dVX//aD99/5Wz/8P3/n3dXmnAF4+IlXOs8yEZgIfCEE+r9Vv5DwFJoITAQmAhOBicBEYCIwEZgI/CERIFhLjsQBAeY9vpB4n5gxySgjYCSCNMjdBagmQnQgblCaw9f4IIi2wSuBeoXmemebQXIFyh3IJtDE9MZUEjdSGiWJFtoY2R0GrN2nfCI7h3Qp6xLQDkMd2KomPqGyskNKwAC3ZDwb2BqMl+6lDfsbTO8C70oA0pZFzsEQ2b3EchBsm+1SpN2wPXyLv+Jnpp1xcUig8odYOsRPCCyCblzJkT6SX7Q3Eeg49LHaJJLq3owrZ+/w8HD15MmT1aNHT3a4DNxKdke+OZnWpTBn22sqMkYdYfSW4IV8XRdm2/rUOiR0FzQoKL1LnShFqPzVtujl/T/nXbLBM6X7XJsKh/wLL9zn65w1Z/rV7Z772PYFf/cr61LZenXnGHKMxl4HZsx5mIVU462zupWvDKYiQGJ/zI9j1JQzGnzoLTFS5B5rh09vumG85Nch5zVz79p3ry7nM33QX3aHj+rDjxqXumq83vul1RxibJaUCU7OGx44zpCH6Nug36ww92LzsE+y/7SLr73WCyVtVaZUeeB9zXtjW/WuCaej1p5t7aftwYm6vs76WdTb/qm5A4v4Oda03RsX9TtGx2Tx3mcHNIJ5sEenZak39XaNLtdUyShXBHLNbQhl5sc92jLtgKkNCTNL69Sea9O2+JTW4c9ijSs//k7QgZ3H/IIsfb7yysvvfvtPvPFbb/7gB393tbl6zF8NNkq8gsm2s4t5KJynicBE4HMRqL8EnysyGycCE4GJwERgIjARmAhMBCYCf2gEjCB3USQcC0HlS8TCLxIYbvcggyjiLclEzjFoQJg35LjzOgHwaK5Asv7nbORot1jfAWtf9z00wbYtwkO+r5vMsJ+Hepsc6zpfo7pdbFsW7Xmor0vLdF3LeO6AWZllvfZjF+RyTrskThE5rds+jY91Leu1bRbruljnvX2W/vT4u93z/shSCkUzsoDWhwerJ+fnq0dnEmQSALxCpq9jhtv+gkPCAa0PkmQxThyMW+0ninLfOrxp3z37KuVW1sZF/31wkYmIDAYl84ZLKsnhFzbV41ijz/6QNyfHx9z7Wh1y8Aq2h8od9jsjSJP2c7x93Wfrb5e8yjl87DbllrLL6+U8Ok4P23OGGGu77b9+1VHz0HP4LJ+E54hXYv0wRcbHGLssfei6tmVbt1tXr90qJQlXz+W+ZJptQ7bOrktmnZ+Qa7RZnqW3+/Xc9rnt2s/rxqN1WG/p+j4re1umdbVM9azfpe6ub3nv7WPpMXqWFGw7O9l6psTXr0v2fDTeynUfV1DrU7c2XH/tX59dh63fvxXwbK7O/eODw9XJ4dGTr9y//7tvff//+s7/9rf/J9LGeO22/mricK1Rdc8yEZgIPB+BuQfZ8zGaEhOBicBEYCIwEZgITAQmAn80CBhhNoPgvmMvcP8CpBUf2KsNqy+v2EkpcahfbXRrbooEgSGfpEUC5EVQrsIRNCtahcDYHJYRVK7HOVk+g7FJ4Dlc0Z6xr1RBBaEGlWTHEAD7pTgDfO/dW0n3ld8nYi0eT7/IQCJLBS0JbKPsKZ8GsYeebcBLeLsHGbPM6tFKtWsQvSOQjj5sc5uCJ/ETraOiZDsDzlfvsgdYt49XMff2yYKToNqogUJ37anFcWf/t/iobwqQWeM4MjZlWo5X+gj89Stf7EOBr9tlDzD1Z2z6cAnvNAixspg+YliBe2VLSQhk/6bhrz4pkrNucLO75k6Hu+jUuK+5o8HuThp+aMfEJn1NcTxEQK4Qi6QFGTdc3axOT4+3dnwt17nRf+e97XtWk8eGhSDhlHUmgxGcHFuc3/aRvNI3/9k/mKJAktPSuksrajIA1USI5C11mknIjG9tpKr8l7Rkv7GM2Vm0Gz+8gIeQ67Xmdp8spi6SMufMjzA5IvtgIGTwfgEE6UZv8Ro+u97F65oPIrbPjm3/4Iiu1zDe6ldRFZAfdzy3VAdPmxhHyKIaFuMrTFCaNd8adue60k8xC0GNrGPbYsrVPv61r/rVpLNZj0r71cyQUWPue2xZ6/piJpnjLdhqnWEn9zR3Ucap8aMGkacheCjL4d8oiyfb/dDA6sAxOydVJ+7Zqy2SVWeWnsYKW/9+OTrtIExWm7q43lyxieB6fbM+Pj5Zn56efnB1uf/33nn48Nf/6r/9b7598+BH6AhpN0YxDMzTRGAi8IUQ2P2V/ELiU2giMBGYCEwEJgITgYnARGAi8GMhkBh10VN25B7/Y9Q9yCDIKkgeWRbKJsC13mP3+lYFk9YpW6HoCDDtY8ic3k/XhQAgTHZz+rZlncF529Cm18ajIcf4smGCYSPd0daybaPrQ2pw0wFz13u27rOKwe9W55AbgTBjLhqn+yvb1/bpYr1lWdf3yvdhndeSPwbRLZOLZ/xoQZ2dQSfeG/pJinG5evDok9XZua941dxFd/ZIqmBe+R6b5Jn3OIBWiZ5dGGI/BEdb+Wjdcry6F/2LcafP6Bc7S5i5Xtq3f4oEi5hzE7valvjkfOf4iPNurygJlrYpObsskpfqz5hCuJRO9fQ86L8b9CtraSz6WhyWrx12e68tbdszftqJ8unrwtFX+UJW4VN/3dI9yZqcc74lcoVdn83482y7JSQSWOpD7GLbeV/OgW3ee16WwmlkQeK8MhaJSZ64rGNpP4id0ifZrH4Gl+d1rJ/+0qNIikHb7jF7/3Rd+SG8y/nRv16zS1+3fXnw1en4W7dyHuIjJsESP5bkmLIeEn+eS541zvPU9+LMn5gcYpx94bjf4jzIzuDT+gZeAY2frZ8Ns698toyfrOT/TdCHEICbmw9Ojo5/42h/7zduHrzz4Wr1BA2wcHt7/HSn1jzPE4GJwPMQmBlkz0Notk8EJgITgYnARGAiMBGYCHxJBJr8qED5Mzqz79jeMYEjaTumNLnBt5k8Rt/8hwjZfZXyVUprrKYQY3Pja3BFZCXIXZAXTVwkYFUPgaSy3hukbgNNlZmrA2FiUGy73kqeGHgqZ9BNJLrtr57Y1R/+SWDZL5oIYnUuXuqkbWaOUGpPIs8SIkUwqN9t0NS3LabZZFyLgDuNu3vtQUmVT2NsnFLEosZXOg2is5+SfmkHmCvzzQ6NS6RiN2NhzMpUHE/b8Mk2jzWv5rn/mJi99dbbq08en60O7tynP1+GxI4ZV2Y5aUFfkmFGP0ko/1n0JbbG2G/fO/ch0NRnX7Ed/SI7IOt+kpMhoZD1FcvW7Tzu84W/ZP7BWvghAQsznHNlh0FokBElm3N0fJA1d5G1yHqEIOKFX8Z6GNIpfcd6cJ6cbInbkK4ODfu61hxIIAcD8eKLrfFNHe5dJlZiaFaRmVkZy/BLGWel2Bl11vgKhcxc6gqGsinVpE+SMpkn7F5f7/N1S7LEtNnqJKewLYNzdHS8uri40O2x5h1S2Qr5Qj91XcZXnxU902fkmE999nVV58oml/s1ssr5HIF49LqvW61L6mm75qFy7Wu39nRDlw7iqISh68R91VzPzssaX68ZRzb5x4570FnKH58nSb69fMlTn6oUWldXzE9k8ZV/8dl1iZxfifT5dwNEx1mJljwjyIe45GMUl4wvbag1K89rR+s5mY+cQ37hq3X6kX/JBNOTIiAd3CV+Nw62ZF27Rh0npYnU3IyfkPg+O+Ll0FCxXpMuSAl5d3PzGHLs//nKC/d+wJ5jj1d7V6TBST0yyFkmAhOBL43AJMi+NGSzw0RgIjARmAhMBCYCE4GJwI+JQEevdidGveE1y2te1rvZN3D0VaREdQadI2g1QLTegNYAk+gzbd4bjxqU+urWMvD02nY5BoNXg/Z0JNhWvoJb2tGLyFN1kmKl1+7a3cmXTe5Hn7zuhbD1bbOCZAQoXed19+1rz3GQ3/ia+50v4zYndaqraIiSkaWoV+p2/ZdjC3G4GGv5BWYCOsZkXfvV5wxeVhD98WuQCPTa+mk8z1t1q/c/+ChYdCTer1MmQ8v58ZU1yExJDjNrJMlQwq2kE3OW+XQeRXQUr50XfbOKn+jTKCWyzm1fc86QUte6aC8RuALJIPpqF53BDDLGa4kXfY4vEFiHZlPpGy64Yg7wI34PWxt4Bz4qwV0VCQvJkPiKfgkLMQtuiNCSrxr6gmPX2VP5IkUKuSKJSm+TJI2IsnQogwvdVVH2WmfbzlphzJI8kszet4+uIeUkEkMgIpfxu75C1uEb7b12zcTyGbpaZJ9JcFnIQcv879E3Ja7W2BxTkWXYG83abT/Et9ezZGCmqAfNX4H9DeQUcydx1r7cMEc9xjLYeJcB9WWszotYDX0hsvHRuiquJX0RH9ZA4zta9b2ebT58kLFX5poKS8Vijrc6+fs1iFzVVH+Xnn+b6gMf1vfebWZi8qakVVu/0Jpr/fHYoDvXjod/9E775eWVWWT4BqHLCr9zdPhwc3X2gFXrAlcmPexg/1kmAhOBL47AJMi+OFZTciIwEZgITAQmAhOBicBE4HMRKBLjc0V2jWzVc+P/FvVrlntmvhjcbZJFNgghCAzCPaoN8jxGAGk8PAJTA0ADcQPRBIOJOQ2UDbp51SoZLRVouheT2U3bgF06DrXUViBqUEognSAb9iP6YqrsGnd2HdUp1nV94tKqjXt971mdTUCoI32wa/DeexYNHoHaKvZpHSFUGFPu6RNiR8mCJfpti17bOSzehx9EViJJ8if2GV9nd+lXZwwpn68gKl8q0OFFza3tsEghkD4553Wu3JsVRIaUBJOtdhx9mRwIl0Wd3SPDaCWgbhWzkZLhpF47oidjynUpdWe6zJG6HOeY+2SuDf231MJtiK42xZAsq8yz5Jljp44sr6zBPfY4p4TYQLevCEpwSVbEN89jcOIowVLrRUfBnb5r6oMxfqX4BUjq1GGxv/de1V0GYlPqq42WIR9dtDkCJWuPuVoL1VZ79e2xsFs2xI/rB3kJZHVlDaFFks+vYHqfevw5hNy5Yt5q7iQPG9ry3ZE4To/Ss1pdoCskYhOArikwaDm6RPbm0rHiO0pCtvnVUIvyAyL3c+uijqsLKbQdBtY57tjmHGzAsHwZZ+YylvipLLWhXBQYq+Rj8IG09W/KmnXAcHCjsKQxNjeslSLOyr5bt8FIpW35Y1/9yLzo28Jf5WpsYMa1snkOXW/9YClEUYd+hehvHzDnSjOtzeehns+SU1aMfU5P75zc3DlZ31w8foDz/r3Ig52FKAGo1zWqmJo/E4GJwHMQmATZcwCazROBicBEYCIwEZgITAQmAj8ZBAgMZVR81ZI4roJ7Q3YixcR0BpYdtHrZGVufIghGgKmMVEFenTJYHsFm1NPmvYeZJp67voP+JomIpvUiwaU6u+z67ELO1tEyy7Nt9rGUXF1XcGvmShEK3W4AH9KCivbT6Bax8rfrCfaj1zb1l9rteNon25Z2c60NR+Z/HOQo2tWvZV33L2JBYqUIj32/gkgG2Q/ffhsl1U/MGkdVlkuZwdKrz2YeDZ9ad2QVdhwLvKq+tCzHaL12urBbOZfgzG9YgRoY7kgvUK+sej1DGFjvdREgEj5lQ/u+YrmR9CtKI3Ox9FNs4svAztdll5gJ51ZGr4Z8Y7rU1dclgzAlujn3+t7KpHXX3vVW27+PGj/9x/qw3nGawSSZYjZWzXOtixCNYLQPOWim2BHyl2b8URyXxGGTNrEpgcYY+zlR1yUb/fu0ascvVdZ4xNe1Vet043ZYzL0EpH1LBh9oF2q07sbgOtje+4w0IYdO1hpUER8FwHPIwL2QR2P+2AT/6bmAHJf4dA7so61FaR8cF8MI9tb1UWus+jSedle+z9ZbnC+LVFm9Ql1EsXWu1O6jTj/64b1atGXxvq/VZR+1dek279M3PkNoMmebq8uDw6O948ePHvJEbs4U4YxY/FRJOWznWSYCE4HnIjAJsudCNAUmAhOBicBEYCIwEZgITAS+GAIV2n22bLcTWFYw6qtC0BaVEWHWB+EjAbcBMCEtMgaB7uFlMOq+Rx2Mto0EqWRYVEBowEo8aFhIMJrI15oKFndnguUi28of2ysgHsF/k2voST2BeAfD2k0dMrEW3a3H1gp8S2fdm2+VIBc9OpfwWbIodioQtj2ZZPjdEa3E2LIo0772dc5qpc1sNEuH51tZzVK2mVlChHyPWbkijGhQBYbNmJFUkdCw+xUyZqSo3T21nhCK/z57kLFZVAi8bT99YFwhLy4LFzoV9rYxpvZdu17nXiFKXTs/gu/KsI/Xpbek6lfqQ0KinMZL7KZoh2rhTtYXlZ75pQdn2t1fLPvb2YH7/UP3HwM5unaKof55JMsviwoTtOuT/rku4+egNMzXMXtMUmlZepy7tVt+SpCGJF0IKysh2cV7S3Rgz1t758CHzOGaeaFe/frjWLNnF5iZedX7kpUOxiqWKnCeGLdzfMOnXj0fDAzhlvgypqQnZ+bdLrHN2VnJuMkarGdhELZ5rors8nVUSzBFXrUXyMe/zBl68dXiOb6N827VqIsUU7NLKf51SCYZuqOHRvfLq0b/ZqAHR0Ok4bjPbP6eiJtYIAscGCx/AwEyybTSEEU/Mo+sBa9TZydt5VS+1vNSffq5c8ElSxTeX9t+7VMdYmgma5UiyGjIbcbBcxYcHTg6XJdmPMa+c+Q/7OfvI8oOIAj7eaXfCX8jX/yTf+oX2Ahw9ZBDdgx/UcaprMTU/JkITAS+AAKTIPsCIE2RicBEYCIwEZgITAQmAhOBP2IEeN/s4ODI7YuIMg1SCQLNcqHCAM+AUKJAEsL71H2GC3l1MBG/AWv1TZA45A0+EzwbOFIMlCVW2o51kgMJUrnuvvYJMUbQaluTZJ4lrwy6lTUotnS/3Cx+tvXDPh5E15ZoGLLto/J9bZPXuddeDbF6jOCZ2twnsEZ2a2/09f52neNRl3otW4zQ1bJ9drx+jTHjx+YNpBh7n6/eee8DBl2EU5T4gz4JjaurC6bVNgT5OEBmOfthSeoUUSIcZSMX6Vv3NQYJHzHO1G4NfMbFID+CDx2KEBv6nS/XgP6oj3Vmyau24kBfXxU8Pd1bPXzErIi/4032Ff4jaHbUgeOw38CsryVbe+2s/RBAfC681IXFlBqb/VtHYR8Zbd7Su5Pfzb9MU8/VUJv7Xpv28SMAPEnMb2WQtR7lvfbLitdX2u5sLjaqd5huhs8+X+qXgFkD5iUyPp8SU1RnLCE/k42Hz3mWaoRFVjrttYYcjvbsGy0STRSTyxxrY2Zd/GZ+rNPvvP4Liey4Li/9LAVEGdfe995h+SgE689sNZ/fSkhVsseFvWFHPLQZxDlbvLMOF+s+1zUPjVn5X+392763vZIpvEtzPU/WezAi1p8+DkIRRfu+5ss5GMhGBifGJgkI3geQbJJqyoTApN2xI8+fyA0rjrnlOUM/HznZe+XwcP0you9xn3eE8THDo46qMUBuZpkITAQ+H4FJkH0+PrN1IjARmAhMBCYCE4GJwETgJ4EAgT6ZF3zX0Tf3oBgI/sKWEdcREBpC02KGTmWhGORJfhjqESam3kDSAJPQNAF4B8YGm+nPr/0qCJY0MCtkECDqoi0B6pDjVLKxYvBagbYEiV/V04Huo05tVCZHZ4dIJDiusccSvjku7aqy/UAzHIp+Gygb8HuUn/rgdd977jo7RAfBtq8GSk5IDg7eITbUK0HV4/KsjhFcVz3kRwgI2iwZCg4OU7GRhrRhCxv6adGb9eHp6uNHN6sHDz6h8zE1RVxsxBa/3E8q9jJoO4CLYxr2xKz8ayIDmXKCC0v51f5YU+PezWXuBWQ31aV/kF+FmxiJLfrEeWTtSWw0rup24EfHRxk/4pnTaxjAZCvhl95oT6CzThe+bu1QdxgyF2n07WNDc5Jnjsf+aMhc4VXs7yEvWRgiMOuy1gFi1U4fcQoh1XWqZzmpb8N6jN6B7Y3PEPVNVKnHos/6uXHTe8hNCbxDssMOIJbM0KQRhZJmeLapff/kbHT4GHkJGvcn8/mKHsfH81BZmNSP9ZsOGhRvZHwN0vlxvBbXZlXUfXzvMWY8tQbdK9DsQTNGJS9v8FPZq2ABweckqRU1IY8gm/yoh3UgwK/4l19uydVz5gy4T53Pc4pm0OnfFV2UpPcimEcfd5z7nr8CGX/qfM4QV3e8EV/XN/ciKMnnc3HNvF6RSZnXIdWttLLBosalLz1Hw+zWpmPq0n6wjvm7WeuTZ/2Y+tf40uhrjOb38e281iSrCgziUyuY54nAROC5CEyC7LkQTYGJwERgIjARmAhMBCYCE4E/AgSMGJeFmPCAdJs9vmRZ7IuBncGnBEq/TmQG2TYwpD0FTcpKBChfJFP1tb3aDJArwLVOueV927JtGURab7BsWfv6YOyUbkkp7zvgLh36NAiPEd0mNkeHNtWtvKV0SVIYGO/IENt2AfIuaLa+S9kqxyRUUECIXMScbZZgN3x5Vj/rlr4EE+q6v+OwSIjJ7rSsJEQTgev9U2DcW3340cPV5QWEgIQUvkSHfkkStA9cS8jc+BU/69WLq8rubFJncQz016e0cb/FSPmSSlv7nSptSnrgdDLE1K8d5kqc1eU+Zarv4gcOau+y8kW77q92RGT0CX46XkvWhR01wU/bbd/FpzByzF0kqWpdZrxUdz/1+fqfpcdZWUjKF2nYssrE9+CxvBb93bqKr6is+REzxkK7w5Uwa1+V01fvDyDH6sMM1Y+Rrvav1+wnBpnDWONTMEAxBBVSyDMHzHWSnSDaskaw4qu3ErVVUc9Gf6nRMXSRws66xbfbz2v7tcPECdS3wsp+IrzDY7d+etx6mYJs9MTOp+eshLbSo5OnslV4uW5qDssmuOFBE48lU13FVW3tm7V55RJcPPffFp+DDZlwzp51+tjjDcTIum6rjtFSmb8jrOPGZ3wNE27brLl6jRMrxxxff/nll7+B6uP2jTNvbNN5lonAROBLITAJsi8F1xSeCEwEJgITgYnARGAiMBH4QyBQka8KiPvOzs5OCOROyQzxi5ZRy5mkD26JDiUCDN4ttndAeT0yPcwasc4w0O6+Fue9R4ptEjOUrve1TfKnom+YTN8ISS3YXzKAxvhEdozaTPhQfh8mxQw29SZwb7lSkD6xP5Tn2i88Sk5I5KBNj7JR/PDVYDf6kFmetd/BseceaGe25auN2jfsRpeBswF74aa/hamBetmzDuvFbkR38IlfegZLpG9g70bosce9eEUOGxbt/ugdX6/EkuQTREaIzEuIpZBSkAmQKFSWD3ZDjhSm9C9cnbDc6tS4oAobaeeMFnS00FZkd9H98gpnyxXR0ULR1zwBupI9hqg2OqNN+y/cf4k26k37SkZUkWRmA5oZpq/q8miySRvqsZ/1vPxWfBL1PY/xY5Chvlbn+uv5oVv5QU0yjtRBe5d8kDDKqRm+i0qyo6jaXqs/90MfEEQLP/qVtaNS1mxeT8QPx+zXGV0bay4u8L2+JGn+EzacV9eJ2VZjXXKBPM+Y6xULkmXr6ARLnpmsES0PAliTKZnDXaZVZYDpf80VcAfTQ22KD6WyVvYAACAASURBVD57uP581K1Lnzz3aHSNccrz53Oof8h4hroLviHj0hnxMpMxq8sxZb649tlz3VtfVFe5rJjEVe9PFn/Qbalr9xUbf28Qdi7xBPlqj6vcuMbMvnPNWJwp51p7Pov6bF91UpP6CPITX8fZ9kNJNl+vhN08OjoK0Un9CU1fx/rX0H4cprf+WKl2lonAROBLIjAJsi8J2BSfCEwEJgITgYnARGAiMBH4sREgaDNa5eD9stPT03sEgXcJ+g4MxitotGkEyISOHSS2xQ5Oc58Alh+K9fnHeVmsbx0VwCdE3YrYZpBaMrf6Gjjzr0vr0oTXZh1JOkhJGRCb8bEsylg8p+9opAv3daNd/Ur7wpfu0/2VKx9BD38tIVsWNjoIV6715axBylN1w27Xe95ADrU8zbmWJLBY39k615j/4Tvv4ggfT3AvJYmJBOW7cdSrjQhKTkkC2I6OzsLxGgoguuva2yZZqvr2b/tvfXElA0R0iUleO43aOB+87NMl5FgNLLYczzVfYcSxlYTDVhSZ2KJltzbUUmup8e/56HE4mrxSqUnJHW1ZxsnLZd94htEQgTZSlv6KR3SEYNJl/drJtX7XT9oYj0Wz6umjCb3as6sw3pGyyvt6KGs9r026F1+tL78YaXKn61ry1a9CujeWerXpk5StzAYu5RlDH+u572tM9Zypuf3q9qwP/cXxJT5SR+oKKadN7Ns3JBhnS8uXja3G4CHhtTf+rmTtMidlu7BUun0tLHv9lu5qc11V9p3yNQfjeW5/8cX6HHS1t8/SFa/p5tVKxuATKGn3dP/S53ylfjB5Xmfs0eXqcH4Z94YvhkKOWfTNOiwdXV9dfPX+/ftfe/3bf/LOm9/7v/VSJzDm01vPPpWzTAQmAl8AgUmQfQGQpshEYCIwEZgITAQmAhOBicASgQqgv2TwRTQn80UQb0YOnw0k5r53c33l19cOKuAjgYf9xwzzzQ4zQ8WA1mLQ2Gf3Jkp9txEyW4wJo8fA0rZkSkme7MgK9fjPkmv1Mhzr3LOn6+3vG0qec42ceyPZx5yT0q9NX3UyE8cgWKpMvf5ilzrl6/U5+ob467FAL8gZ0blttG37GPh7fqqM8RoyRy/N5bcjpxBgL+slBcxy6YwdRSRwIst1ZBfj668varbHLLKOt8semWWG3L/35ptMJeQY+tYHR4wVssSd+y1kjyUDUAzBJpk+ZpSVYs5mnNUYksXluLrN/l7nTF9wcLy5tZ7DjDXPRcJVnfMe1syMJye0OtSZ38bZMe/vH8JfsWG6WT1OHntv3bl7ul3Ojl3ysXRinTG7NBovlWb+8Sx4DgyTV8VrinlF0bn2nxigy7LZ84ugVaeH0iAZT3xy7hrnsW7QEX+HDten9/nnmaP1m/HVxfp8CIH5EbqQSKzla7CxbxOpWKwu6FfGV0yvY8Nnr9qCBdjazlSXTX0f9g7Vh9/xy+xFdLliQkjFj+qb/sOckMdvRD3HP3odQNKlfvSLt1zrr3OhnHbqudaJsls2nXdmYCEn1sEKHCvrshzYZ4vD2ASPnMGmSs17TUvVuT6V8W9Ry+zHbuHqnNWqL1tC6p5j/j1gKWC3MHO+s55UIpAUXyG1znFqo8aRptQHU8dLcb0qI5HpZv8yzuu9Qz8u4UaNL9+9f+/Vv/Ff/817/81/9V+u/sO/9ldX12dP6OXTG8uqoI8HP9vxpnb+TAQmAgsE6ulcVMzLicBEYCIwEZgITAQmAhOBicDnI2BIWGHh58s9o9W0KzYC/0f/7D9++MJLL79AIH+fIJHKvQ0BINwH25JREgjf6t4BYweSLdNBdYt3e993P89LWe8N5C1d3zKto+tbl0HqUr7rW14OsIu6nlVaR5/bZt9vddG5r5Xp9tZrWx+xY+A7gt/uZ33LR2b8dD/PaadfbAyXvW6Zrte+WTwG2u+9/zE8JxvbQ2fabvYWDkZ77+/V/UMMyBRIDw2f7RMb3cczdRbJLARzHxmvR0mbcoMM7PqceywL+fRHXKIjpBFtGzam35J+47VP14FLYQ9Ww9fqLL5qq78SLY299b1mIkO7Mtp5Xumxh/CRSVkUMWodLWezdrt+Ib7F0bq23zqCtw29FjClnshRXYQT+8Lhs3Vd3JfMDzy4R5mk6uHhYcZqnf39UIVj9/qQOq997e/4cJ3DLDyyQpONZx/7W3d8fIhc6atXA6vv8rpt6FNsoVvfal7W8etT19lLrdacY2icPPfRmHjfuDTh5n1ft/xSTp36IFnasxUMubek/yDB/cpp7iFb4cxi3/t8iXL4k3H5fw5QvLZde8s5sM37rjMHzNd+3bvOOvzlFFzoeY1r4LVevfjo7MmrX/nqay/+S//yX1zde+EllTjrqnu6ID/LRGAi8NkI1BP62e2zZSIwEZgITAQmAhOBicBEYCLwpRAwgDNw+3QhpYtskH/hX/3XV//8v/iXjnk97wUCyPsJUok3kScyJNAkESX91x08msVh0FhkTGfzqD8BpkEiXXONbQkcg08vrRs8QQgP07aoTukgddzSXjpim0r3G2udntfJrjGorQB2m8GEbIWj9MeYdi31JTt5CggX6wx2OcwCscMVWSEG/ZJL+mIRu/ar68zm8dpA2fb2v76Eh5/m3PUgo6XHTyAd+d18ZN9udaGz5ykakfP1x2y6znV8QadyZoM5Zq8lMp6QnPLOux+Al+OQQCh7tW8Z9xdXNVzkt8XxSQjkH7VbPEpG3ckupGnbywy1iG5r4gNgwPKwXPQz/Uqd9xkT52SmLcjK9kPeYDtu5dGFW6sX7t4Lt+laTLt+oDt7WeGFs2O9pdYWZNL+Ua7zJpv1g8RwLSgbXO0w1lVe96M+r6VSfT1e3fP14siX+hoj7fEDH7TXa8I6utHGERDVXzIt75wzlUNIpYVfZTKKm2TOaM6y2xGAmW8x5XF0XTWJs8MiHWjXbOmtubO+2g4GCSRRZBGPJVeTTLmBSbdHlB+fB7/a6WuUBxByzofPtgSUu5gVWeXg6pmocYjf02tavdnzT7wU8j7kp3NpFhZO4W4yGcWH/4hfCdbpU7/iypjz/Df2zgXflLTeV1CjlAciHxlp3PUb1eLg+s+znAla2BzGbFOPy1sf+8MgNofz4pGTvJQfpioD4+uj7Mq2fpkBv/ibv/nb+w8+/EhGDSVOECJKWvpcd/N3IjAReAYCkyB7BiizaiIwEZgITAQmAhOBicBE4CeCAOzE/upXf+2f4JW2+y+dnV18hYiXjaUlf67NILMkkEtgvnXBwHtHAnR1B7QSBQaofb+8blnP6lRG3mSEwts+ths/LnV0RFlBsdlmlfXRxJiyttGpzqO/9VuiZfgVudFO5Nqqy2/HTFHG8XdA33W7VyQr2G9iRPn2wfH0dcaJr12WtoPvaFDeQzSWupb91HVAhpBivjIqyfLkbLX66MFj4nGyriBDpBxq3zhGRnYWylpFnb0fpCIeV/ttGSW3dcjo2/Cr/U+7jihnu9ccUZ++ZTf7nNk2dEpKpEBcSFbuB5taCyEnEZX4s0vhUyRZyEteDV1k74x2zdYcq7dINNwqK9vfrd/tCy3WhTjKEJq8KfxbPkTI0HJ7LVjtyJSFFEGXBEitg5rLWueOo/VJLlsyNskbSJP+wEVkFv61Dsfuq5Otx/omvNC01d02PDt+ySNf1e36rEX6xgN1DF+jS2aV4tqxdB9JKzP8nJuQjdvno+a8pPt5Vket9fiI/i6N3XIM3aatvPorGz/88t5rj2eV9k8yTt3ee7S8M+Lak8j2+XeMpRsP45Z+Vj91MOJt/6Xd1tv2kkU2XAqB6Myv1/DvYDTq8eelo6Pjrz98+PDVm6urd/KwOgjHEkbyU8vT1lkmAhOBWwjs/pvzVsO8nQhMBCYCE4GJwERgIjARmAj8OAhUPPb0/8wkmIMAOzAaXf3BW28eXFxffZX9sV7xC28WXstjO7KbG/fvMbOq9usa0R/tpbOC6G0waeZN2kpHB63qs3SAWXcSBP5/w+UXYWral8FoX6tHG9mk3OhUEsKDYr1yy7P1IR+8oHS7wWzXt8+xoQ6OfTJlzCqy2P6sQN669NUNZCLHqCUOzKjxS4f8Rsfyx3aL9rq0X22rgnTtSkZA2lFs66Jr7b/nffJUfF3ugtfILvxiJWSZmT2VQoYd59L+HFrNWM2U0QeOtu+1M7e1ZT8PO3UZ11sZ64dvy7GhdadnvBoZFcNmXsnsvqkrv9QriWHRr+YTe+7L9yIsGwPASMqObenHUCVB1GM/51PuM23IuD8bKyn6o49761zLy6Pld2N1zkkVotT8m8mIIYp6sr9VbO9ImsYmQqwIp6XHkDrWr+sk+qCfrpiXPAOZiVA7EbM9JAz4+JXLHJCH1rtHmDpYBjmoEhJMSx5LjCHP2a9s5vVUiS43/vcZ8qCox2fphldbWy77wfm08dx7XLEZfWPsq5wH4znShnoaJ4lLfbK+SEXGiP4c4NfjaLvpl3UGSYqPG8hPcTJTS3zN3Npw7kPi10Ns9d56M7vELdiN+e2/OxJjHpfsERYZ9XEUy6ff3DME/ejxed3j6frgogYwCtHGnLvvYsMoxrwu7NJOV39YZ/fPLq5+7vj07s8geApTjQInmUZMisEsE4GJwPMR4ImfZSIwEZgITAQmAhOBicBEYCLwE0NgBGe8hyR9wB5jBH1fJUD8OhkiLxhIWpqs6GAxlQanHNsA1EBxBJepuxX2GRgv+y+vmyzw3PWen3WdIB7LtmnH4nUHtR14Lwmwlml96ui+UcBP9+9z13tW9rb8sn15rY2QAGO8rc+zx9LX7tf13nffZVvvAWWdfrQuZYnrZQdS7/3DR5+szrMRf+GtbBdq4M2YN6J5ibdkV+2ao9e61q+vy2Mf0qHLbRnrlU1pm0NX6rx2vlrGSuT02ZKeC3wkbpT3cO8seJiMtV9l1b5k1OUg0qID3a2v/ev7GOHHekuda/3s7qu+ZawX756z7fhG/6Wcst1u/bZtYND3/Uy1TNd3f/2FzmJstb7ljNjNyuatTu149Nhun21Tr/XCK/lTfazzqeXsWlCHZ9VLYHJ43Rvyp37YTQaXTlDMc+uMLu+14/PW69R77S/9qOdyPN9DsXIto57ysdZQt3m2tM7GrZ8Dl5RHl273C5VeO9omsjy3Dc+WzkD0uuv6uu+XfdTZfwvEztJ/c1oeXyHIynGm0a9l3ue5+zbHtxjInXSqHwdXShaV83IiMBF4NgLzFctn4zJrJwITgYnARGAiMBGYCEwEfmwEFtGkwRnZHAR9FYFfXR2/+dZbX6XutZu9q2P3XyJdbMVrQWxpVe9aGbwrPuLLZE4Y4UU0wWOpck+hJGhUfIueERxjsvsnoCSCVJcZGBUrVmDfQajhI3SDPyntqnsVVSkCw+u08TXC9NFvbC4Da6+3eod8y5Qugl3pAwgJfVO+x9nt9q/6GkfqA0D7XX5s+zF++9wIxigZd9ug2mwxv2hZAfawrSxKrLd/ZZSlinFxz9iuyIiRzIhPeC5B8aO3f7h67HuW61P68IqlZBkJK/m6HhlAhu1u1H9zSSaQ5JJkhfjzTz1l1rGJX26rTjupKP96HnKmnlnMPAVv8UDfUwtAM3nl0yakg+1YCxEvuiGZPAObNRvJX92cr45PTuL3mpSpqwsJinJMWxa3c6okQlYKy2I5p4Vpkbxei4OEBrMSvK1TPq9+Dl3d33O+2DqIFe8t1SeXXFed0PXrkpmv2AgKwpuSep8fF4d7Y1GbuvEMxFcHYrYbRZIsWYiMU9N4zBlyivte/drPegBT/ZPysvQ6RlnVY1P96ecP+mIv7fao/pVFpV+Fo/lPGcCmyCz51WAV3LjGvsNhSWYpOYuuk2SnOfDr8kcLjldZfwpDfOO+XtfkYtnGtbocazBKR20XQSXs6rN/JB07Mn6NtOZpEIw265MZZHagl3LN9SrrP8lfTbQ9JS2RpUE5CbZLniWP3pvuwGw4MRm4K283D9eZffik5SljeOOTTz55gwf61J37JbUZ2j718cpOs0wEJgKfj8Dur8nny83WicBEYCIwEZgITAQmAhOBicCPi4DRquGcYd3pz//8t79xeXn5dV6nPFahwSmBHnt+EwobTC6ONmhdB5LWeU2YGtKsZTx3375enkdguZXxvgmQblO+r9XV/fs6FYufZbBrv7a/lL9tY9nm2JfFtrbf9a3Te9vU57mP7mP9ss1r2zx3X7oF71Two30P5doXr7tsfZFwovOde4erd97/oF4d0w8OCY+wR6NfE5m3s7la73bE7ZtOeajGM/Ut6/VoGCeICOY99cu29Csd1QGRxdisU6eEna/WNSYZM3394mJtnwYpyIV+NH5e29d7r+Mj+hq3EBTDlnW2W2efEB4ShcPXltUfry2Ne+u1ruW9trTerle27ffZthxC+DQUVT98CCmtTh7GvFqIz5KkTZT27Otd29OH5bX3+tBHY9NyIaMh4vwqqDLJokKxci3bfbftyGmj8WhdtltvP4tniaHW02flvL59H/0LecnTrKFo241LGx49d/rh4SuYPW99bj/Ubem+ubn1Y0alPvlcFHHqMz7W+pDt/p4t0eurqPyVM9Ox57jHB1GtYTlsUTXp8fTs7OxnfvFP/YM/+6d/6R+7VwRo1gigMeBZJgITgS+EwCTIvhBMU2giMBGYCEwEJgITgYnARODTCPg/JZ/1PyerfgSPBmdEiGS1qODw6Pi11177xvXl1TdoODHgvCJbgm2t9jowNmjvPZjsEsJlZK8o3+WIrxwmEDcTCaGQAiMW1PYy2OwA1L4GmVUMPCuAHxUJTPOVQPNgzLTh8KuD5sWoc4ypxEcA2wG5lbZ3ELuUX/br8bRs+7n1QaBI+sieRiNg7jY3QWKzNgDdEYZriEcA3vq3tGtArj0Ps48ah2v2ebq+vtTQ6hCZYwiik6PD1dEBWWLgY+RtBk2yaLgW9wOyqxBdffDhhzIC0cVXSEOSrcksS06L+I+2+Mx16nMzqLGI8CNLQKm5dg4Zm/KpqzZlGjvnt9u5ilx+IGEABf7VPthAB71KBJ3eWzImBsBOdxB8kFYQZcmyKenV9cWOtJIkcz26UpJ9ZDqQmUycJJLMKPPs65euVw9HZ/2NRDCZbGVakkIdHkrQpDxr3koJux5TkyDb8Q6/bc8aizdxI/MSZeob61k5+7p3lUfba/3KxwbQSL04txb7tKyvlLpYmgjyq6bJHqOPch4mJ/lcSN54+Ay6R1YfVUtlMqrsT43PUh7WwkB7kmf1ZdgigKCQWHtOV60t9tnCkP6YZcea5NpMKg/36Vr7XPLsxycw8JVMD0s9kz6z9dxat50nVA74R10BkTmkzT6ZLyy6Z5wlGDFaR23Rx2DJuYt79OXw+dEXfeLIeLi3rorX6nVevVa/Ootc5cKbiNq/yUD3Hsv4WcPosqh7QxrZtTeXl9dffeNb3/ra3/ib//3df+vf/ffpX36Uzfq1zywTgYnAZyNQT/xnt8+WicBEYCIwEZgITAQmAhOBicCPhYCBoaEsURxxq1H1evVr/9SfP3nta9/4Jm2vE2CeGoi7Ib+CBILJIPPGksASHdsgk2sDvA7yOkC13dL19ksAXgHktq31dT960Ofp/zmsjKVlvG+91nvdur23tL32s2pLtvW1Hvt33VLO625rfZFbvB3lvUfsDD326cN6j+U+TW2jz+kLqUEG3+rBgwerDz74YHVx9oR+sJVHx8mkMiD3UK/Fs/0kfeDRVt/97nczraMx7dBTpseEXDFTMPLW3dYx8E0912LZpV+J9N5xxn7L97mF1W1Z6N8SbNQFO/voN6fcI16vfFa7OG1YfzhBva+1oi4klMRCkTI1jloPPe/6pb7W6RqWLOt73epxNdHkfde1HuW6tL7Wbb22gwHX3d7yy/P4vkL0L3V33z6jkf/4HJZe6z1adzb/Z1zq4IMZYFPjuA29Y7LY96AJpHpsUm9/D0ufG5u2hSfp3z5EWPlxYb2l+43qnGzreemzDda3G0u7Xm/1obbbPKu/56h9a/3dp8/aaH+saz1dt2x/6pp51M/lfC59Ulcf+iJxrc7dxwcq86zH2nbtgxxLmBL2eP/o8mr16uXVzb1f/nO/wjRDWudV2kZ157/+zTIRmAh8GoG5B9mnMZk1E4GJwERgIjARmAhMBCYCXwiBXeD1tPioDykG50BqBnuMrf65v/xXVv/sX/iLdyDLXiew+wZfQDwhWWXjflzc719DsNwQwK+9N2tEwsVCsLjcvL0q69eg0YDRs31SRlZJR8t74eiKWEpg2u1xrYgOg03tJOgkTM+9WWSo7IDUzBoDVzOEkrFGm3J2tdgWP5ThsETfqO/70p3mp37ajrGuSsdo4lf0iQv1hNpDb+F8W5/+lN1S3xlA3sV/fYMQevL4k9Xbb7+VPcbWh0er11792uqEzeqPTo5XR0dHcClHY+zYAd+TO3dWHz1Yrd5664fBRX3J0PEC0k2fa7MkSE9tkO5CWiDjYCz4zkSXDJlBDtGxxE8zhbgekCUjTY0SXpJmZiClDAH3zOqijBxsbFNZ48ai/bQiRGQuhQilLkZcJ9jz1bmDw2PIoMvV6d07qwvMZH3Er6CMuNli+JHh8PVHvt5pNl4X5Xvrt5p7SZeYLLIHX+kREuYazEM+0t9rZxJT+Kp/YMG9Xz00C8kihlnffT1SvsKF0GZW4zYDMkSIDxN9Bz7RmNvxjNDfuqwBzjqYL0yKlBiO9X25ch85Np6HRC2iVNJMyBjY8EUdUKjbNeprhE1QWp8CztloP3BTV0Q40+HzUSJmm4l01ovEKjh4LebWW+IvdZlb1NAbZ8qfzBdifk3VbDJlldOWKy+y6JB4ctpjh/tlhuT++nDbb9uOjn6W24fMEfUhQ1Fm9lu8gSRUn4UrvUuxv6Wz2niLPOvLJdl/2+IrPRxHbxVWdpSq50M1Hq7hGhvXrJHxN/KGr2bG5DVjPrpZv8g83n/rrbeRgc1eXaKc0ywTgYnAF0JgEmRfCKYpNBGYCEwEJgITgYnARGAi8KURqKCxokiCu1/6pT+z+sY3f+br737w4Ru83fY1g2MCQ14PSuZY9iBrGxU41p3XHbha0/fbYJg6r5cB7VMyBvfK8K/1tr7ledlfO7dLgnF8UUeCXMa07N+67df+WOehbvt3221Z61u2dbas5xTGWOQI5AG2LW3H69ZZhFjZlRio17jwGfsZI2G8Qf677767evjxg9X5xZPV8dEpm9NDjfi6K33+9D/yD69eeuHl6HQa3XT/4Ohk9eCTi9U7b/9otXfyFTCt12bjrwSNzjFWfrg2oq8MHcm4qo/D/Eh8FunVY935zhhr3ez6IJ0ysOxbz/bLAksfbady6BCDwkidknWpkLijk9ljviIoWVFzX90jm7mtTCjbZFeuIG2a/FFmibP3EjLRyXXeJkSdWWprSN9eO766KXkTnTp+q5TeqnRsWTMOYpSMd/RTVkqGEe4w8y711cFLpYJvCCRunCp9ZIylutaKN9aXDXXWfcg82iR4Snf50+tJS91veS0hmnFauSjxhXvRx3KRmdiNr/zkNc8hX/bqJrzfGLs19AiWyQL0XgUU58H/RGLUeaddj56LjEIibTyX3a6spf1cXmujx+r8W/TDjwb4anJ8os5xL/srpx372ta+1rl0et2H8l4XQVl+qy944ri6DvwgBTJimH7W3+zdOz48eu2TTx7f3z84fMjb2DxorpHyVb2zTAQmAp+NgE/LLBOBicBEYCIwEZgITAQmAhOBL4yAgWWCy1s9btW3CJHZvruer773ve+9BBnz83R7XeLGoI44j9iSC0peFZNYoRgMtkyCvxJJH/ebIlbfBd8QMcuNrO2fPsaGTdLYfxwai8FhR1sey0BZHRIifSRryAwQRqVuZW0zyPe+daTNujF6673u19dst3iWnNE/SwfPyXQZgbR1ORDL627DVjrwY7CcYFu2BzzahzV7s3HHvQRNvSoZP7TJoa733ntv9dFHH0X/y6+8svrm619f3b97uvq517+Z1yzfe+d99tdyD6jSm4yyw5PV2++8u7o+I7MIk+rM/mycvY5BV8YY4/ZsW8bUMojkkh8LujpJzNvo8mKUnW5V7/BDKRLO/QhptGPBVg6pEhVbb8aWPtPfr3IGOwyHKEOeD0bE3eDZ/qNKcsjXLy364evAPUfUYGYx/+iX0HDOLgE5WOsLRb0hy2jv8WWp6wAlU+geU2zCZXsf1Vbki9dZN1sMtOHrna6vGnvwwSf1+Yw4qMKMcfR6o07pDXuxVdsOV/1s/4TVsZidJWl6yft7yXISS2xYur99vPasDkvX9fo3Y084sv9XWDqIopG1Zt8+AsnQrx6fsjxpzgVy+tSynlPQ4wgLBjFfHvpTPinbYzTrzZLx4nPr2vbU2UUx4zF7zA1fxdyjfbrCZ5DBB32pEjyocw81S+6dG+q89nAI4uprzxKojsFjfzy7WTshM2uO1cUstT4uyP9jLHvI80CesC/g648ePyFLd48UsgMeACceKc2n1/yZCEwEPguB3V+Kz5KY9ROBicBEYCIwEZgITAQmAhOBL4+AsRjHvgwGsev+6SuvfuVbFxcXv0AQ+KrqBgGWfcc6OPVcQePTmRbKt8zta++7GDxb1OG1537FKaH0Z4SI6u7Avu3Y18Ni3fLoujSOn9v9+r7PLdv3rdt6bS/rvV4ey76OsGW7bwf9PQZ1t4zXjYV14v6R70rC0ByRFXbIa4Z379zPa5UG6Pfu3l09evSIVzDPQuxFN6SbG5b/4PffjCv7h2avOL2DJBhY25jXG50HsctByMG5xrsMP5yfIjiarEDp1m91NQYMwNsU63p8fbahr8tOyW6vsd+6HKP1hbncQWF/DK/YbVlHI9OrM8ys82istZB9zEZ9WUQbRIWHZFrb9Nx9Oyso8k0mQXAoY+k5zM3ip8fSOqup8GzfFuIZ5LJ3TQAAIABJREFUS9+37r73rL6lTudiOx+0tUxnkvUYJIUlh7332uK1utqO5yZ6nLo6NqsLsHf9+XEHfZY49hx5+3D05vzORddrQwJMWUvXxzrruOekx6NMj89zt/dc9hzE54Xf9rO0/uV1Y9x6lbF47zro4n2XlvG+65+lW0wstvUYvddv93lrm973MfTQxP89gCtXEJAQsydkkf0sq/TnDo4O7yyYZxfKzjGVzzIRmAh8CoHdk/ypplkxEZgITAQmAhOBicBEYCIwEXg+AgZvCdaeEoUdkD3Z2/fzgrIGd+/fe/HblxfX3yKf4vTy8jx9iO38qJ+ROtFh0smgKyoIJMXFBgJGXxPcZbZUYIixPYLKEfJZ541yFoNMs5uM0m3x2BBoWurFwFzmxyDfPZgM+jMWrn1lSp3ed1Hn8n7fFCAUb8xgW8h1xhGUW7q6N5Jy/UqePsZf6x1hiUV2aXOrE+Li2i9XjuB4vcV7kBJk1hQ+ZUNFtd9R4VBZTliin4dfXnx8dp6MlZPje6vz88vV2dkFWUfXq6M7J6uPP/549eDho9WrX/366pD9yO5Qd8DZvbZ+9zts0M9+ZcEyGTiODYwYhFOQbC5xhEAjLUujwZ4FQHuRACWor3SwBI/Rpk4v6dfZdVHgPTr0Xz2NU3SMKcp+ZMol+wjdEi9ZD9qhnnntPa42ki/gkMwbqBcz5EjuWp0cH60eXz2hq5hDxtCnptGV6FhZm8xHkxg5I1PjFvd1SB8Mli3O273xBhLiaHFPKe0cDnLMOZT+yf5YGW/EgLfmzGXi+DtrqVp3a88PJcgf7ZneB7Y+RxbXsrZMf9R09un3HGyUEFewGjhC72V8aqg1XzJXvBcdIggfxE2Y8/rlyJpTCuvY9sx882+TrC+novz0XMsFm0jFN6WzBor8KhX4rN6sEf1Am2PDtuo9Z0zc9PMjjiXv3ltDNmMHM3od3vDkq8+Jtt2sM/2hLvOGr9U/A8BP9mHj0vaSa51F6mk/+jJSv8ipXvtWvX9T5H+Da7D1OeXCecautqKbWfdfskxpplf86UxHx6p//h1UXsx77mjL/8EQfeq8Xp88ujr/+vHpyTcuzh+fMEMfO1aKb/3q3CwTgYnA5yAwCbLPAWc2TQQmAhOBicBEYCIwEZgIfD4CBm/PKhW4Eent84oPgeiv/ZN//s4v/OI/9C3itG9B9pzWK2HpuybogwOQ+NjFb17f1qyMgWCIBM6W7tN+9P3SJ9sMkC3RwXW/IuZ99zWLowPP2KfN0jqV6/qu6/Zu87719XBuy3pfhIDExW7cFaRXZs1SjzISE63H886GunY6WncHzOrpUv1H8I0+9imKzpdefHH1+PFjXpvcrM6fnK2+Dwl2cHIKcXYO3ozH4JzZcM5+jwyyPfYr856GXcQdrKgj+N/f1AbvsTtASFZZsmTCcghqjtTLtFgkD6wP47GQq9YtVkvMRlPhOYgJ60JY5QJs9C02JBAww3iiY+wNtuIjAWLPG264AMElcZbxlHaxLFUSMLJ3RdS1H+4xZulN6r1O/zGstAWHqtBWz2Gtt7EOsJlsR2S7fde3dFq/ewZK323idcPz1tyX4w2uzhR99av9Vk/8jL9askgYgRfFtlqnhYcfZBCKG4hp6a/WcwER6nXIoOF7FGQ+vCo/sya5Dqn2lG2eazEfNiWeKput/ChdeOZtxiDeuemm2NeO/rplfXyPTIlY7zNvfc1m1cdvLvWtng9NNAHaz9VurDUv1bdw6rna2XE+DphjX4WkVWeGf6Vvu3fZsHPNJLnmet3FV/r4zHtdVGKRr9pv/8Y6QqmcKv7D5p1fnx8fsgcZMq8yqKPyKr9Pg7lomJcTgYnADoFJkO2wmFcTgYnARGAiMBGYCEwEJgJfAIEKd0vQYO1ZhSwfAjKiOwK/f/qf+Qurv/Kv/Rt32eT9jfOr659jb6s79HM7Hz9IuH/IZtMJ1hG3uHl49EqYULZfLbQDgSOhJEE6wTDZPEpYZzEYNWhUl6VIMfqE0CgSIw38GGxXN/z3P+hu4qJlemzq93qbCcK1xcwxbRnE5l5FlCYYaIxveX3QDBj99Tx2cG+9NESudVnfY1B3+5GAW1nNDH86mI5/Q09fq6NtdJ1jNlvqq197jc32f7h68OBBSJmr8yM26j/Iq5WO4Zvf/GZljrEnlhlnB0D68OOHqw95NXOPVzJXB8d5jTAEjEo9xDHQg4f3KXXuMaQKPwPVVobavubstDuFGaeC1DlkamPAGc24cq/dQWggV/WIioW5gj1pw51wb2Bq9k7mG83MYLLm2GKNVwCLALuC9IFpoEVVzp36dEUbXFCKmMzFkKlXNNVrUa76Vr99iDT7U1vtgBVyzUxCqmKLgetbxhEsWQvIQX9EVzriSWUF7ohW7ZiB1GSK+Dl0E/K06P2azDJ17UFgWmrZli9KqcNzv5KsUzXWIvQcVmSSKYU8hIxdtFvjqnHudNWzkcxBnPA59F1A9zNTzz7PffplnJpWqP3ZrfvWbeak/kdf/HUQjo6CPmam/o0qn/HlM7OJ34gChvZ9PmrMu2vrtu4g0+2Zj+Fa1WnS8Y15Y9nsHTSG+OODAV4OCS3I6qS4K9N4We/fkJEVRhuiELj7WZshx3z+xz9Tbe0P+0Y/128w2gN/CDKeUxhe6o8Yw8t8cOMV3rE9HA5o3M6zTAQmAs9BYBJkzwFoNk8EJgITgYnARGAiMBGYCPzYCCQs/DN/9s+t7r7wytfOzs7eIGB8bbMxM4kXz3wHiXiQvYZI+KmA2EC0D4PVLgaEKttmBo2GDla9jUxFoqMV5eg1Y8VNsbeFzdBbtoPv1lOB8CAobumyf/oR0Fpu+2n8Wnoq66OkfA1tZCQ5BmXGuCQC9Y+a6Gofonzo97p96vqW63oD7KVct6u7MbSuryXsXnvttdW9X/7l1eMHD9lr7JPVDYTQE7LITk7urH7hH/hFNu1/fXXv3r2BH/4zFY/ILnvIsbfmFbbgCtFRaT06SZ0EhTYhBxioBMhNXt0LMCUzmEklhTe+ylpxk1fWQlDUGigihJEp6InjqfnHRjAIUVY46kfjkrmHgOipF3ezx8TBtsakz0DA2Kh3KLRHT88V94cQZiqTAGMvvbSrS/LKovzTh8RUrWHrW0Z73vfrnnZvf7rNduc18LZuzuprXepTvovX3rlZfNY7RCxLD90lU9elQ3utq/W17aVOdSvX/imrtvTlwrP4xvYYl32U8ygbA8vhnzh2fWT9ocQPwVehBPiYo/an/fN5SluJpe9S1r3fuvAi7fiiKD5Q798C+7e/nvWlz63H/rdfjdUv5VyJNb5as1pzTcR/VoOkXF2r5dPFtrZnq9epG3rVJUb990ESzQKiOTeBqt/xnWr+hm4uNhBk15uD48ODF994442XfvlXf+341//W/0hH+mOCzrUQomX+TAQmAs9CYBJkz0Jl1k0EJgITgYnARGAiMBGYCDwXgWUQWIFjunQgdk07yV97q7OLsxcIQf8EmQ7fPB9faoMd23BPPFokkVkohJUJ+IznW3cFj8OVEViaUdbB4togWhLG4JvA1Kwx93CySFNRkU2uF/7FxtC4vdaewWaVp8k6iQpVVnKLwW3ZczOnDHaEncahhrHGocb58Um/Rlzq2TF2hpHkhxkxawN35HpvsWjBn06m0bdhwiawySn60zbGq70O8J8aL73xeNuPgcbWV15+efWVF19KlpHyZ48ery7Y62zNq12H7MW1NqWKEjLo9Gb1yeMn+Trj/voEEob5OjgM4bAn4WjCIDiZ/bIZyYObME746xzhwWpjSk2NxF/nMH5KqIFB+Uyt43VMAOR4/NpiCnXBElllnirj3n7J2IMEcS0UIYYu2jujbN+Jwv94oj9kjTn3F8OMui/MxkHHxdnZanN5vXr//fdJmjtavfPOe6sXXnghXwD96P0PVr/yq7+yYnO9Wju45GtxIdn0P2YlS3aeOh5Nxk/XpyULnkqKtl0LCJR/VU0fyC7xpb+vhEpEXimXPjkhA25chlAZdtQTuhYbeBY/88zwqmj2xsNe+vAbTLk3M1L/JHosjqcz7vKMhLApYsl2s/SUj6WQnUVAuV9b1vqwgXmnOUUbtOZaIlTbTAFnvImMawb7uUa3Y2UMIbewAU0YAkl/ghnZbD5+fW8d/xm2vGBMzKftkmS9n5cC/u2J/5rWThdkxdv5kMzsttLtDOgevtGW5xcb2aONeZKUuhkZa4yM/gfYHeOgn69Vaqp8KfvirL0QbKrAQP2tYejOOx1qTWt5tbpkwYKHGWRmed7kNWzGCHKnr//sz9356//xf3H81/69f2f1n/71/yDyAw48nmUiMBH4LAQmQfZZyMz6icBEYCIwEZgITAQmAhOB5yJgYGnwlgC2pDsOI6Y2ylsdn5ycvsEG+N++vL55RWIFZsXIcJs1ZjcDV19B67LQlyqDUuuW9Qat9pMgs31Z6r7qetP8ECcItS7l+7r1lg2/cliZRst2g33tEammn6RB94suw2Xq7KNc+uKC1EwXg1kj+cbs/2vvbJosOa4yXH373u7p0YxmhCxZxiaQw16w8hcLVoSXBGyIIGDBEjZs+HsELACvvHDwDxzADuNwyJKFrNF03/7ged6T596antFYcniZOapbVZknzzn5ZlaHz+tTWa2/+1jvdY7uNM5dnwwt6rwve4Wf/q39aV+K6MhcHNoPcjAWG75Q6ZcDHz15M0SIPjr+vUQCY/UVyzfYmP9Xv/4F7frHNu7OOe3c+F/pZexFJmKLa8dZjcNXiTDxkyXhNb/4IB4UtA7xgZX9KYcsstzVj+Ouog6uIFWChThTkQw9ZbI2HF/PG8347Cuu+q/Na8eADr+YCM8XQqexkRD51YcfLv/2r/8uEbH81d/8dXx+552v5lXUf/qXf17e+/rvL9//4+/FHbE6rhGH+cJzcZxzXRY3/4Xr6Hn8vLNDKZ/znNC31kDjYD9xLMx6HfQ4dM4N5EEGu7W+Ij8wFota10pSUNtrK3Nl1cBcna4nqKbg6r2+aTNQqnPobe/aj9aZDC/E+r51a7peiT0+Q1lnQ5/tsQPRJAOtz2V/nHU8RRx8Ntvv43NqH/2t5cE6l5xkJUhWux4s6rQ9uIgp+Fj00/r22/b2vUSqf/0ZY07Sq35cPyVrFhvPAUU7XmdOhw3H10fbahKts2DtU/3Annn3Wl2fffZZ1vAb5+f8aTzZXu7vtn/4/rexFP/X7sT+/JkITAReRmASZC9jMmsmAhOBicBEYCIwEZgITAS+AAIGZZYXgmviRwIyI8WKAm9PLj76+JM/IDHpG4TRDwiraTLo5N8Ne+cQsBpsGxQaQHpUgFpn6yVJrDOwzit2aFbODdNLtoJNM4PKpyIm0F5BacWtCuku1q1oOwb4kgsGzqVXGQkj7ytAr6EY18YPuqvBPagMTs1MsiglAVEbuXODPTy2KcW+BuGSE+uguMYAkbMKuGOHXo4zRVwS2HvfOsf4qOm+rct+QXqM+ZR9i26upXDMQpGM3CyX++tlyxjsk+wTW1F9utlhqzCQ9Njwutfu/GL55NnlAq1p7/TxC4XOh4QDjuoEngxiUC+ZuyhSb/wIoIhkAoMNawLBIuL6FUtMFHGE3uqHMvWJAXo8Chf0pQxi0HpfkdQWsn5Js+QlJ6jXRXwSe4kY3c78wo48vODDA1kehY3rzvX09ttvLe+9997yne9/b/k6ZNjDhxe8hvpg+eEP/3T50Y9+tFzyqqUryjnVpyIuuEaXxK368+VCpfSLkq8buja9jZzEj2Ored2ip5+pWnnIufY9cRZvR86IqKsMJ7Q65Njo7KjTEJ+FUcaMwCk+qdOp0j872Zb1krWgfOEMmPHPrK7gSIu4OF8nZgNS4vOmnpWaE6Y3JCr+YESy1X3WDmPHnuPOaFgHZhy6qb7tWC07tiPns9I4SGA5QY1nSKGasGQzxr+hJ/OctagddQ8CDfnyUTtiUGvF+fDDnyWLDX3kUI9koLazdyA47cDUfsl0i/3ySSzsY73tKeCQcXMWyMKAM/okZrMcsO2fwuMcoFumNl2cB7r6nKH7Gt2eb8hovE4GWgi2u5vrLJyTG7IeT892ztEVx34H7n6RtpTogf/NMhGYCLwOgUmQvQ6d2TYRmAhMBCYCE4GJwERgIvBlESC6q2CRUNHLi29+81vfYAPpr7NNzrnZR3zmUDbJLIcKJkcAboTaga4dLQaOTTD03jv2sxisK9+v4FUAmqaXfuzT7UaJrQP1qa/Mmgpiu+3YpwLeDtbpnD5mHSnTwe1Bvtx7wZ4OWa0Pul/nElzba10dvNvPoryB+6tK91dmrVdZ9TTRcMLrfyEV5UBSCLD1h0PCoYgTpRkTc7JlM36zoHwH09dXnz2/DKl2clYEQm0hN4iBkCvgIomhn5IPsKKAwz3GqEt0rj2vh6+6sb6XVLmDnEy5F87bp0tfp29XjrPrwvFIqAR06qWU1lmB4nIDQSiBp3u+RrpjqPZTpzpq1mljHI8fP47MDfs8Xd/Ycrc85RVV58tDf4TVlhAkIU+OY4s9dO8g7XCM4ziXRUBRRV36cqX91KA7r/iNod8fNzOuKwcM7aNM63Es6u1+7s/vfDO9KWl37rjrtWdD9evzELaevj7XqlWnclkjjKkI3HomrVefpfW2D6m0Hk01yq4p7JTLYTV6ypcaU7W1X9VPzF27Zlj5dq+ku/+66Ou6qK90lh6vMyrXeTQN/RBb7WPWg3+6WDc9X9bpT/QlE62utRWdq3mRmHVtqc8+FsnDQ398UHfpH8/XmLe8Vkm7cEr2qccxSpJBjtU9TKU4X5xf+KrlJXsDXp2fn9+6rkc5TmLXzPNEYCLwEgKTIHsJklkxEZgITAQmAhOBicBEYCLwOgQ63nxNxOVLbKhA8mRLnHb+NYK3r1HxIMEdASL3JEooY0DLDwHgzdiLKESNQavBJ03sV6YYImSbkAXVWRpyEBVslh5lKuAcZ8NRnSTwDLmGVx2QVpZNk1tmcBTBEZ8zMOwbkarTYSSUL5+Moctu3Oa6MoU66DbzJu267TggfLx376ewRYxDGspiQJzsofh6DLBta31ty+DaMuA4ZOY0gdh7mEmo2OdWfO0iAYk55TbsRGWk7TyEnNA/2txHSRSdixvSaSqjDMIAUm2PDne9Ot0+wH033i8cVL0h2+z2+qpet0RvESiDBJAZQ/ktthBAmkJfnBuXXFPcGyp1mR8rUj0Q4nrYi8P2rWkJlgecrQ8TB/GlvtHHUWVmW4eqwdx+riNSGEMaPn/+LASEpIfExdX+ajnLfDF+MnbMlHL/PMevjHOze3Cx8FXWHg7ZeK5PSVPM1xCiP/MINmyeXnYlpLDv63HOfyZAtzjSb7T7fPi1VufJ/cZcow4zj8sYg3rMwrIkk4+z9nyVGZqFLC7HWIDqlySKMJG8ydmMN9qpiI/qipAQFUbqdd1oRwySfahMGjxTrw7qSFIs/bhTr4CWjn4V13WmXtd+MsvAkVevo9v+qg0unGMCmxJ5GWMqhl8Sr7YFMWT1H+XaMflKUZ/34yvb+Ijn25HJ5nOoPdexRYyaDr2FQbQNEUw4bvUNOa9dnGlXwDUtfoV/YSbBOr7Ki1b7ut9az3HpPJKqtjtGffWZ89oJdp5sy9jRz9AyV9Zfjz3zXOdN0juGhw8uTvhC7S16bjiu4c7uTv2gBqV15Wb+TAQmAp+LQD3Nn9s8GyYCE4GJwERgIjARmAhMBCYCXwoBo0kOT7vlj37wJxfvvvveVwnmvnp9fXVOgEfMl935iduNBo+ZYLnhp4M52z0MCvusTF8bHK6Lcl3WOqzzfn1WRxev+7Cu9bdMfanx5Xrttc1XXeufR8sY0HqoV3/6WPvhdUiTUals37c/Ntm3X7NSv219DglBUO3ZYffYh0oq6pVWiZ7OgolfBuEE/OpRt6++cYKAMfPsZPnw4/9jI3v8gQmJLwPTMkJnfJDsa/8kDmKb+q4z+rev9Z6bhIzAkMu1P76i5sn6Uutg0mz/PnCYOvdFKwJKP7IBfST5sY8i1muXOcictD0Ih3M+OOCttho/Mfnkk0+Wd9/+yvLTn/50efTwjXxdUB3i9vjxG3nd0jm2n/IW26Mjd8ef2OS25ZWzLj61L7Srp+skybyW/LRop9u81451HpZ1W9ev28QU7S/0aTk6R4c+eXS/9jGNTUqt/JHY0Q/LOMWPkq9fdVhaZ5NV1ulzn/s6FfwcfBsV6tGWci3rvctOP9Tr3Ow4tsGOjr4SOuSV7SP9advSt0n36NgeZfKMoMd5WPfr6x67ci4ydepzn71WVr9pPYwnaIXwPM7bGOJhTaQP/SQTXROuG8+SmmTkcn+cp4x5t8NcbJOj6+ChAlnXzMoB97YxzxOBicCrEZgZZK/GZdZOBCYCE4GJwERgIjARmAh8DgIV0n1OI7EmLRyb5S//9u+Wv/+Hfzzn+vf2d3dvGfARv8lqET+S90G6inUGfhVgHgNotRtk9rmDzlfdq8OiTB+tTx3uJ2aQavE+mUNmQiVDpEajDjNRUiRm1Ek6h1k+kgqVndOBb4mVLoLe0c1aA9hDhtXwx3qH4tcq0ydZM/pbPulzsoWEDXckpZQzsLfYXhfIJ8UEGYWQz95MnMuF0r9B3kygZLZxztjo13pO6GSbast29Tabx/2itO04YMbQU2PWnQ8++oix6XMRRMTp5aOKxBfZa7MAqRY/9cRzOw9bNKXc8apiHDAN0B7Ry3i9d4zpW+PHiaoTaNuxZy9/gpPkBNe9DvwIRLKD9Etd9uM/S3yynpI59nVOMpJ+/rP/hXRwrBAr2Nuwz9gpcv/9n/+1vPno8fLjH/94+cF3v+OyTrm8vFy+/53vLk+fPg2GZlFJlqi5PgQAqQIm2nO9lW+1/5l7g1ny5UPaxTpu0ttXW9tGhguOPa7K5HKosYIG57HGor7j2CQqJTFTiz7ngblhzfgcpI/4Aq9ZbxovPaxzdPazcpANeGLY67HWGYhjExvMOfRR1kBlpCGncU5ptz+32tDHWo/Yp1o4JWVTry7aNy4s+1fntK3H6fXRN3y3n89WLvxqbeEirr7SavZdsEFMvcnk1FTqIdR0IrbARj3gVL5WP7vZ376dTefg8pzbxtFjU9aa3JPVRUvIZQd64iPL+lWX/kvgiQWa6h9205acQfshzo8y+bvC+OpsnXaKFPRvAPruYMPY9o8nmLQx1iIJkJvTN954HLn4mKv5MxGYCLwOAf8czDIRmAhMBCYCE4GJwERgIjAR+N0iQDD3Z3/+F8s7X33vARkQT1G+NWjkuCUINHI8BJVNZlmXQHS0NTHQZ9vVsT6v26y3v4f1fXifgHUEpv0VRrmBHRvQ29YBd/dpO23L+257wUdCW4tt2RMI1sEgtmW7nyRgZw6Z6WRpXzs7SB9adwT4Weuxzmw29V8TOEuwePg6nXbMNJH4ihz31nnU+AsD7y1rO9W35LSnnkORMOA1LbmHn/3Pz+0Ye73vW+Sok0TMV0IHSSHr0LZ9NVYFjq/k0a8fumJfD9kUS6770nrLkJcxsCATW7n0vb6Ws+l4vdbV/XzdUxlfrTyV0IoflZEjrhYxkOTS3/fff385v3jA5vwPl5/85D+WX/3yo+z79Omnny5vf+Wt5YLN/UOIoaczfBpjdbU/6/O63es+XD8W75sI8V4/Gjv12N73tlviM/VVjkRK67Ze8qfvlbdIznjd/W3v0rLruhfb1liXPjMIfZ6DMb7q57p/29Fu1/eY2l73fdHW0S91KmPx+lWHZKXPtm1uVq88rFERh752yp+gzv5Sj+36LafV+nM/9Ntufcv22XqPvl/LOJ4eb481RB7y/XpnOvLTY++5cP4lG+uoddHry3MX5aU1HQv+ojZzbCrZGddbM81mmQhMBL44AjOD7ItjNSUnAhOBicBEYCIwEZgITAS+KAJEms/3n5G9ccXGVZs3DNQur/cEk6d3pxzZzJ2A834AaVCaoI+2dYBpfRczvyS5Ouj0K5dVDGANVjtgraBauQpkKyg3c6P6QiRASmx5pUqbC/sPIbHc8IKS2UW9p5OhfzaOh6BRTwf3Ej83fmFu8D6bA8EBiQQBsxlkkaSVAWxYJnTZv7KIBjnCfQXWsVRi9DG5SRtyFmbZbKjTb199tBiXV0YL5Bz3Zj5RMZKssEHoLM4pNEmm1etmhd3YMjzjdFw4GD/cv8lijbif8Eol23Atv/jlB4Uj7b4+efhKovIclXUneYX+VRAfrNXfrnDN5kghqdI25k8fSgeG1Vc8KoDpieOts1lsmiwP0xD59OnqErBTtUUM37Kuer3QTDbXHa+hPX3n7ZBS+/2lGlIkKSTHvvntby2Pnz4JGXZzs18+++x55vOMfmYf7ZNKZ+ZSETeuouz75Xjww6ws3ekvhmbMWHA0AxLmrfxk1qkf4+wxsI6yPm3BRhKTWCpYy1oKLozLfaqyuuhXWKqdtcd9SB/OitgLBytDCVPKeoSoZb24Pr1HJcXrftbKLyae2lrfLEmItx6FGWVkZOk/+nnxlHGrWz1OQ8mpvzOpkj0GfvqnrOV26CMnKn0ylvQtP5sEPpBR6rZj1ovrBry9zZ+MXC07cLMyX1Z1hGJhRhwmt4OwVkVeacV+9mJTh7qG357bZtfZ7mGxrg5RVrUOiHPZ0xPx0mYXsXCjfYtq1JXnMjbH3yU69N9Jz2LmP0k+qb8z/rawFjFthuCZfwO2PLcQZMuWPcmiuyzkcv5MBCYCr0FgEmSvAWc2TQQmAhOBicBEYCIwEZgIfFkEEt0aKUI47A3sHhL3kkVmwJ2MHTgQA+nKclkHmFoywLSuz14r322e13VpGHXGlParYJvA1PiXIPJYpzThZ6JFM0+MJaUzSoa4nz5FZrQP0U8AK0fTr2BejywkA/VsBj78ra/4HQNc/VGPRR80awZYj6f1dbtn2wzw1UvonX4JiFXmfxCeW6CyAAAXfklEQVQpaUNGzYWlYy1qxXPv7yTfoH1npN5aw4dAWQRRfFIvxesuh+tD28ny/Pl++fjjTyKnDV+/7IyrkE5SdBgsQg/92qF/7A096Wd1CK8iDUpQP4cPXjDQ4N8OjXP8GmNybE6kBIMlPqRvbo912D7B14w1fhfp4mt2N5J4+sY6MBPs9KyyCfVTok51jufswWZ572tfi7x6xroOeWg2jwSIBKg+B+/hR5Mp2kg9NhuD9lJ9LZfxdQNn74NDk5yjrutb1AxCi2SpgznMS/xw7KyNjIe1EMH6KdK11qWEntRcWpwfFs1IqMOH2rOu/VNXPWNHotF+8RWSRpLMa972w25UZiz3/Q45NmyW7rJvD+/bXl+rs9vKfuHT9bbFh6Gm+3e79z4LPkP2P46j9NRrzq6nuldfF3W0nnVdX7etPluv/tzjT17nBguhzWuT2JCcd66KRKxnXfmMgbN+WKxT16uKsmbKSUputltes8z6TgYZ8rs8H+JRql6lYtZNBCYCKwQmQbYCY15OBCYCE4GJwERgIjARmAj8Nggk7O6OhmKJ5sgAOeUVocfEd2eHoJ0cDZs74OyAsIPPY3BoIFlyHQx3UNt93FvM6763bwWS+lNESOLMEYTrYOzgIXEkspUhBaWQzBH2vKadAHX0daN3XzdMfImiG/bNchxQayPgRFYG6KbIKvUb/AqAdkPfxFYF42Y+3ZJFx4tfIVTM+jKA9WuTRW6oAb/VYX9tH8bklwwJot2YO/r9hbigrzLuu+QrehI1yRSj1T3PJNNuDNQTmJe+jAEA9LoxLaz5qqDZPGOj/cZWmQ8/+Gi5fPbZstk9QnMVXy3U9jGDT59x3HlLlpHXokcRbGTZeI7LIlbEmsqQUbW3mWNKVfx9Kainrzoy3/YLIVRdHF/m1ltJgvHPzKz4pNp0p4Uxmj2EKirxAV/fffddSMDndJXouoodcarxMc/0NdNQXaenD4bOIop22eAf3AaeumC/7q8ZMcyXJcWA+17brb99XJ/N3vO+v/QotJbMJWujfIHVHQ33dUoGt/70M8XMeUfPhi+Vto9+mVOC8Yp5Oe7PxerIlAXYrKnAJWiwTD57FnXUZOWWezAaVbHDD0insdda95PUuU0Gpog4FbVOe5zWOUZcQ++wpZwYUim+jZeyXeLTuLE9fiCf/d2ozxcvecbIZM01XsRDXxu2rzCLva/jts9tp3XnLHE51pfPWQr9fS1S+T7MJHPN+1q0z7vFrLErxm43Ccj4WSlvy4Znxr8jbCuWeozQw3713GTvMv82UKOfyU7lmW3f+EAB/7FI+WowdaaxsRD6geBulonAROBzEZgE2edCMxsmAhOBicBEYCIwEZgITAS+BALGa0ZxxXJw9Qff+MbT68urpwR/Z2wbvdxdEiCSPgQZlC9YdpDbgV3b8t6A0XZLBY8GjYNAGYLdr8/KHYuyLxNABqMSQ+qqjDbuCXINNB1AZXiMQN14VDWnpevktr7WVxlQRXLYLiFQRb0E1fifzf0561v7XcPhHr3sSJa2zYYgf+yR5Hh7rI2BeltHkw8oH3Jl1T43sAAG1r7uJ1l2QnC93quoX7V8gUQBg9gb+vZkQ+lDv1KXV0/FkH+//vWzEBLbc0gbZPjwY/xq/wp7carifXDwFn9QzKA7e4862kOKsUF+2iN2JLPsdijISuCoo+y40JhrWSuL+ilpQyZ31kFwMLG0058xmBVmdp5jFAf3pNpfXUIWbZa33mI/sbPz5bn+UEJu6SOHJbhpkv7Og6XPXqtzWM61/VxTFq/tJx6tT/n7pdtaPtlpK6Gu76r1Gum6V51bTlzUkVlyzzguHIp1vYG/HBrOJtPK8dDEeMr/1q08vQ7jtF4b90vX+bx1aV9edR+ktYd886qlo2xl/WNbfb2O9cXjYEuMh3LrUs/6zjX1LdttNZaqX8+J+ul0eHaV775pQ5ejaj+6LpliwWf8fUDmhjWVfQKHPp9/dbVtCbVeDl2nL/E9Phe+qrWuiVcz9Npnzg6b7szv7e2G4yH3b1xd8Yr7snxqG8csE4GJwG9AYBJkvwGg2TwRmAhMBCYCE4GJwERgInAfgQ7uE2rT2OfUwxcln+L0wfnFE0ioJwRt25u9hFBeQ0vc14GgJEJfe14Holrte9s8OnCsPgaRxyD1mIVV/vSrZerhg27RFVJjhIr9dcsmvBJwYuNmZFARqRNskp0FmWC8zAtRIXWydxE679iby3YYI4PSHCFyyuDB38628Wt/bL5FNg5EEf0cy43ZI9hJoJsYtwiCjNsIPOOmH0VioHHwXnUSY8qiJdlkd0Tf7t3lvkr6ZFuplTg4ZtzYZoSvPjHx65W3ZKd5LzGjP8r4lUPrPvjgA7JeroCkfGGTI2a5CAgDdpTEV8d/R+B+YpaWbAvkBAqqzblWdtjOmPLabdVJXmWU+HPYi8wacI6fjDJm8DVF4AZGabAS3RJ4uR8ZOVYnyy1rQL8rs8r943ZnF8v2dA9B9oSuzDDrVIIm67I3ewO5WlsaY370jzFpxhK3cz7Oj7g77uA/BNObeuvsXzpenQmV9qHDa4tzHFzG2rE2TcpRSrzmk5ZhQ4JGEhhpBCRuK4uvnhH3+VLWtaWcY3f9OP9FtA679DNbsfaw07LkUZG8rtisJ4hmPZF4Uxar8UEN5WKt+R57j6vxoGuKurTvnAXHaEXvyJpS2bqvnUq+xqwXvX7Tf+wxyLAyduVTH4Ywvf1Jsd4x9GvMjhRjafNH39p/iS5LZ3pab+aXWafBo5oPmWM+r8kw5blRpV+Tzd+U9HPN1TjGshI9hPSl7PqnxkKCGBX1LPervRGs5pBxfDr4AbYe3d1cP0SNBJkTzvCCnZqOgxr95mkiMBEgU3iCMBGYCEwEJgITgYnARGAiMBH4HSAwwrdD4EUUtzzlNbynMBZe00DASwRO4NayCTZH0Jag1WtLnzsQ9txBbwSGTLdbV9cVXHeA2rptk8hJppiBPqVt5Iafta5ub5ntdpAmQ4+y/UqjgbJyTfY5Tr4nl0wxR2p9Cn1EwSESQyeItt81RINjI3qPmCRF7I57K30dMVlpXueeX/WgU+LEYBuewp5YJ0DnVU5oL9rFw/60xH716bGmnrYO/PUttiG59D3kFzqePXvG3FXGymET9NFP+egzo0ViBPm1/gPxFWIM2RghG09yUJ/2gKGTo6ROGUp0269uIn+wp8iQS7u6MtjcVZuQqxq5Wj9WcIuv7mqvLQ9JQcknXy+9xp+8mXZSe0SFqADjJlmjgB/76YuHRQy1cb/etq67f+19r+u1TF7HpK3nRbnDa3zMsddZ45KR/LPY33LAJ3fjXohZwxbnVJvKeS1B6rWaspZ6PIjbQ1m0M2/IIqWdqivSue/zOvLoW74csdGu7mlHv9dn2yz9lU2JrB5LtVQ/x9l9tb+W8brvPbecdtwzMM+mROHwL/aRW993f2067uA7rq3r+6Otow/5AinP4J5sscKm5F25kmLiKhFfvh19laCs132rzb6OM37hn69H27/t09M/oHmWfR1Wucaiz44VX80ce8TZTDL/AIXOW49RnbNMBCYCLyIwCbIX8Zh3E4GJwERgIjARmAhMBCYCvxGBQVi8LGdcSVgXsmPHnk5PLt48eUK20c59c55dPaeZHY94tc1ArQPJvl4Hqx2Mrus0dyCbYqgCx8TvBI4W1A7d3g1iiiv1dHAol+Q12zCltH3P5GWkTt/0Ye2jsbX62Qw7bbu78H5FrtBQPgsBWUGQRCe7CuiTZUatPigTX0a2GBptSQAN6xHbEkj5twdHSSRU6kft2RVFkVOPR4Jzalq3cvFfpoG+tY8aF4dpKzvOUnxi1CcQQ7rUGDnQXEPSGcRf83pk/KZe3XuzjQjErYN/qDau9SFBPNdakYgyc6b1JStoZI05DxkzGWI9dmpcIjk58GDBOMovMRg+5qLElNOXFe86Gjg5YXGksDITTF366fj9cqOUxM4MOucGjK6uiuTw1dusZNp9gfIGDBz7NQNyY3R9U7UEhjjUHNU5DmDHeottB2xTY50XypQV7ySsasz6qUx9DEFUO2PJiRQ7dUaIfrZjYYxNn9Yb65cf7rHnglAyYx2+bZn4musiQJvgtC5ff7SXA5XMid4i1nxFucauG2rFKbBQ1CKhZtUBRZvFeNj13NfpEHHHXQu18VzLZMwRXmE65tSvxurHWt77ZL7hV8+BiYV62ZmAqtOvLvbxsKR++On6qjbrba8sLsnU7F+I32qxj8dQoZrgZ1/3NUuWJbL+rXGN+U/f8hXU3NFBWY4aC9dgVwQb4/b5Zr2b8Xo6SM/D2PBVO6g7wwfJMYkyF1ieQs6zTAQmAq9BYBJkrwFnNk0EJgITgYnARGAiMBGYCHxhBAjhXig7snKeQGg9odavqlVAzw1BX2QNIr3soNd7S98PscgkuLwnfwwKj2RW69QCJlPs+yo7VCaYVMh+IWy4VtY+lvvX7ZPERe83dM4m7fa/gXHTJ0kO/0d2qKJhO8QH1zU2iTdfN6SPRJqmCJSL9bhvG9phEBhrX6IHfdpNdszwt/yuAP/w6pcGtM24vLSP/XssjrPHG6xiT0z5QiOyZp7pvx8TMGj3NcmTk/rio/I1JnQ4YkkRbMRXcQx5JFa1t1dsoRMeoIoZUJINEHSxTZ/IoBclue5xexbTQ+E+bSErEGdMKRIm2pBsoE6/JKHc6ynOqcM+6hMLQJHwkhwzk0ydVaiwP+M9ZCHpF0U8nDPHrt+Fw9FfZdQTn7HRON0f4/q++2ghmI7XVJURr7YVYgXd1udodwc27b5js71fk+366JNOY+2p0486iJzyBx8wiXaIH21cs8YwUs2IOOdFPgd/9HTpMZeNrq2zbdp70U6TQGgtaA+d1jpyTf+yV+NuwbWc7euS+cWmRbnqf/S3ZVuH89o2WlfBUn3v+24/n+F+vttO6Rvra6wRJzHZXcMPB6wND3GRsLP4nFok09Tjod2+dl6cDAlK/88G+x19rnlkHe9ud7cX9JMgc7L2HBaVe9xD26ZZJgITgUmQzTUwEZgITAQmAhOBicBEYCLwu0JgRKcGoLdb9np6k7jvTUiKrds5GdAR5GWDfg12wN+BqAGgpYPU3PBjfQeRXptJM+Jz6iuAtL02ux4umM/CZff1bJzsmd5RfT2+WmeGlP0laqIfgsh7cjT4amQFzAla6dr6yjdDVSqxU5lt5X++KieVg62yJ/8jSXQMiHONHV+v0ps9wXDwgHQxIyztymsIx/XHEr/IHkmho1/arD3Oaly2y/3cQq6ASI3LjJnYliwq3O0vMaJWX8/UtljaPzwS/mzNUOEwvD6/uABzM+bQgbx7J7m5PaNMhk6IA/RhKEf7K1FVnmvRotOSaMjZoA/Y1D/Xh6V85Tw63jp2bHVmnfb9Z3tkzR6TxVDOQwAorTdf1IwdSSHtneK764jXKhmHfSXGdufny/bsjLm4TF+0R75sdN9hFzNMX2yVzsIwhvmxLs36RdFGy4m7mWsBgObe084BhWui3SyuxlB/Mz710E3S0fsen0SdBVRT3BTetqITIbkKDocTH9BS/kl4okvy60bMsC8ZmtVl5iJrwi9+IkD23O1yTkakJfaRQ0kImvZDPzPuQZj5BEU+v4qXhy3PiiuM0GNdVhPXaI6e0S0n9SKecfffjcbT+S67Yy3d699twUk9B/9KX9GDdIoemg9/U8oPu8QmWKQrePd8il9ywRQScefb+ch4wNN55t5TPau0I2v9TrzSNuTQkA85HPx3fmp9+rfJvxMqUpd/Y+rvjL6BY9aL8pW9ttnsdvh8QRZvMshqbsCfvgFYXbNMBCYCLyEwCbKXIJkVE4GJwERgIjARmAhMBCYCvwUChl4eXc6Iqt+C7HrLbAYzdPiimm3wZRXIJeilooP97phgecikAxFhB7nH4NiWI4lge72qpgtHMsJ6+6gzX5g06DeWpSR45Vx9i+C4NdPJCNR6KIcO8tvH+30iyE9efzzorWBZWXWvM7yUl1iJzV110K+8sgf7oZ3I48LgExzNwde2rx6vJROPmJQ92yw9LnVaJF2UtdjW7Vs+ntDXtqlXmwb2ISvtD2lQfQtLsZagqs39i9BDwMnkYH5DPkIABEv8lxyFuDnSOFqi6Ie2pEcydcwD5/hsXw8nLHp6TDUGuzcenmOrZb33mpJsstHf+8jip+PxwwMPzs0AhKTcSygWqVOY1Tqyv2SE7kXn0K12dalHebFKhhDXseHYVocy1kuQSRVJknmf4at7ED2p4155MelXMMv2ccyH8Q0bbdOzR40BPU0IUWefmHQwoyhnvYSVxX2vygdAYWzueWW5giQzm9FXAfNlS+rKh8JZmb5vX6yLwZzKvjI50qiJ8fdgQIH3o6XG2rp6rbe/6zGqL+SSuoct5dRtm9dHHGs8NMRO4yNBZulXGx22IuKlbdtDypL5GbmBi/rLlzq3/cM4VEBRztLj8azOEz4i0EUJ5bRnhmraq9uhn2Oyr69Xti77tx/W7W9viPNvL6hLBlnbRqycscMsE4GJwEsITILsJUhmxURgIjARmAhMBCYCE4GJwG+JwAi+DPjYEvzk9M0HZxdPlrtnecXSII2DeLsiUe/XAazMSAI+AlADWov3HQR67iA5hFQk6sc2QsRxVD9JF/XzX/R1htKJ2THa5ouS7UO0UG9Q6+bX1nv43t0dWVpdUqcV20Zp/6RWtJevBsYfBTqrpsZqjRyMr0WpVT0hxzhLxjk+/zn+m2GWfCe7BYfCpbCJe9ipnB/7FxGAYPmHgPr61UMJpBpT+Zn4GzsE0yF2tGPG2OX1ZREBsDMh6/D34cMHEDi8cnmzj767zZnOcy+JeJw3N74XD/9JVYjHLVl4Sb2hnqpDyauVyjlBDiYDEvcaa3QMUsJOZo7REkKh14fjER1mySaBtfPQp7j3RXop23MVtPWTrLiqO1kur26X55f4SnriBlIpJIXjQ85rS9brWJtm/Tl31mlaGf0KxtzvRmZbE6TZeB9dji8yZgJ6M0BhqaV/kWIQXDCk5lWZHdQ6xcyxeh8CJb2rveoK83pVVN1CoHecJWMcS6r1o+aKFupBUd+UQVZdyY5yPCHEyg8zN50uIdj6dUjk+lnchNEtmzGIpxbXtbho20PdXGWNHXxLve32qH5YQlZfRl8M9xg9SxDZxvLNHBRvpYLj34/MG2vCtcgnSlWOjXrO2pc1vtVe830gS/0bwD99Vo39nHuz7eKPY9HRUbJGxn3WP508J0svBhwPFzyAWTsC6i2HK0ldwcX1MPQUTs496wr5Xnf2T0fqGSuPepHbZOttWMFntyfXZ1HW7vUZ+VkmAhOBlxGYBNnLmMyaicBEYCIwEZgITAQmAhOBL49AQttDN9mxR28+IFA/p27TQR+BXl6xNODz6MDZft53SWC5IhtW/RGREKiguAPTbu/+dd93Jetd2SjbJzJEo5gZY6lgues/P5pc+9pkjT7HbnTR9+74P7UTyKK/+lVgLXHlfRMoboJusU6dHSw3EaKcAb+vqhVux8Bau2Y6BbdVUG19l6OfEkYE2/bhkKyzzWwwtMef7I2GH/v9ftle8Dm8R4+wvV9O5cXSW9IL+8i4l5ol/ooBulCcOqkFZfKao0wGmEs89J5kjvXgIdcWfzOe9n3Up3G0pR/tOUPq1Ouedu65a2mqMOBUdx99E3tolGW7M3sOvyQGL/e83goO+gcp4iu218n1Kl3tU6/NPqtXLDf0RVMViArn6jC31PYaqLlzjvWpxmAWoQSluvA24y9FNU9et/0AVI357frqy9Oh4moZ7YNgomPPa+ZFn8VhyLd/ve4kP1O3gtQpFLcel33lJFPwvTHWJ0vf54Yf69tPRrkap3pL3vlal5YXz75WT384ItmM3A+TdC0F7cPtWJ9i3XXqb33tk+c+1nbWfewnOZY+XCsXUjHzVvfK3C+RHzJIjeaRfYjdtufz160+3b5e3D6Jj6Sg2CvffTwzD3aDa675vNzfnCB7upOlzeofJuvUJl6onDcTgYnAsvw/x5QWhN97J+gAAAAASUVORK5CYII="/>
</defs>
</svg>
